--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2012 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_8f54fdb6bda2d271.vhd when simulating
-- the core, addsb_11_0_8f54fdb6bda2d271. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_8f54fdb6bda2d271 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(16 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(16 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(16 DOWNTO 0)
  );
END addsb_11_0_8f54fdb6bda2d271;

ARCHITECTURE addsb_11_0_8f54fdb6bda2d271_a OF addsb_11_0_8f54fdb6bda2d271 IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_8f54fdb6bda2d271
  PORT (
    a : IN STD_LOGIC_VECTOR(16 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(16 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(16 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_8f54fdb6bda2d271 USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 1,
      c_a_width => 17,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 1,
      c_b_value => "00000000000000000",
      c_b_width => 17,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 0,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 0,
      c_out_width => 17,
      c_sclr_overrides_sset => 0,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_8f54fdb6bda2d271
  PORT MAP (
    a => a,
    b => b,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_8f54fdb6bda2d271_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2012 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_e7514e290b172ea1.vhd when simulating
-- the core, cntr_11_0_e7514e290b172ea1. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_e7514e290b172ea1 IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END cntr_11_0_e7514e290b172ea1;

ARCHITECTURE cntr_11_0_e7514e290b172ea1_a OF cntr_11_0_e7514e290b172ea1 IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_e7514e290b172ea1
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_e7514e290b172ea1 USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 8,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_e7514e290b172ea1
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_e7514e290b172ea1_a;
--------------------------------------------------------------------------------
-- Copyright (c) 1995-2011 Xilinx, Inc.  All rights reserved.
--------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version: O.61xd
--  \   \         Application: netgen
--  /   /         Filename: dv_gn_v3_0_6a34997a8a73ba6e.vhd
-- /___/   /\     Timestamp: Mon Jul 23 19:46:28 2012
-- \   \  /  \ 
--  \___\/\___\
--             
-- Command	: -intstyle ise -w -sim -ofmt vhdl ./tmp/_cg/dv_gn_v3_0_6a34997a8a73ba6e.ngc ./tmp/_cg/dv_gn_v3_0_6a34997a8a73ba6e.vhd 
-- Device	: 6vcx75tff484-2
-- Input file	: ./tmp/_cg/dv_gn_v3_0_6a34997a8a73ba6e.ngc
-- Output file	: ./tmp/_cg/dv_gn_v3_0_6a34997a8a73ba6e.vhd
-- # of Entities	: 1
-- Design Name	: dv_gn_v3_0_6a34997a8a73ba6e
-- Xilinx	: c:\xilinx\13.2\ise_ds\ise\
--             
-- Purpose:    
--     This VHDL netlist is a verification model and uses simulation 
--     primitives which may not represent the true implementation of the 
--     device, however the netlist is functionally correct and should not 
--     be modified. This file cannot be synthesized and should only be used 
--     with supported simulation tools.
--             
-- Reference:  
--     Command Line Tools User Guide, Chapter 23
--     Synthesis and Simulation Design Guide, Chapter 6
--             
--------------------------------------------------------------------------------


-- synthesis translate_off
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;
use UNISIM.VPKG.ALL;

entity dv_gn_v3_0_6a34997a8a73ba6e is
  port (
    ce : in STD_LOGIC := 'X'; 
    rfd : out STD_LOGIC; 
    clk : in STD_LOGIC := 'X'; 
    dividend : in STD_LOGIC_VECTOR ( 15 downto 0 ); 
    quotient : out STD_LOGIC_VECTOR ( 15 downto 0 ); 
    divisor : in STD_LOGIC_VECTOR ( 15 downto 0 ); 
    fractional : out STD_LOGIC_VECTOR ( 15 downto 0 ) 
  );
end dv_gn_v3_0_6a34997a8a73ba6e;

architecture STRUCTURE of dv_gn_v3_0_6a34997a8a73ba6e is
  signal NlwRenamedSig_OI_rfd : STD_LOGIC; 
  signal blk00000003_sig00000706 : STD_LOGIC; 
  signal blk00000003_sig00000705 : STD_LOGIC; 
  signal blk00000003_sig00000704 : STD_LOGIC; 
  signal blk00000003_sig00000703 : STD_LOGIC; 
  signal blk00000003_sig00000702 : STD_LOGIC; 
  signal blk00000003_sig00000701 : STD_LOGIC; 
  signal blk00000003_sig00000700 : STD_LOGIC; 
  signal blk00000003_sig000006ff : STD_LOGIC; 
  signal blk00000003_sig000006fe : STD_LOGIC; 
  signal blk00000003_sig000006fd : STD_LOGIC; 
  signal blk00000003_sig000006fc : STD_LOGIC; 
  signal blk00000003_sig000006fb : STD_LOGIC; 
  signal blk00000003_sig000006fa : STD_LOGIC; 
  signal blk00000003_sig000006f9 : STD_LOGIC; 
  signal blk00000003_sig000006f8 : STD_LOGIC; 
  signal blk00000003_sig000006f7 : STD_LOGIC; 
  signal blk00000003_sig000006f6 : STD_LOGIC; 
  signal blk00000003_sig000006f5 : STD_LOGIC; 
  signal blk00000003_sig000006f4 : STD_LOGIC; 
  signal blk00000003_sig000006f3 : STD_LOGIC; 
  signal blk00000003_sig000006f2 : STD_LOGIC; 
  signal blk00000003_sig000006f1 : STD_LOGIC; 
  signal blk00000003_sig000006f0 : STD_LOGIC; 
  signal blk00000003_sig000006ef : STD_LOGIC; 
  signal blk00000003_sig000006ee : STD_LOGIC; 
  signal blk00000003_sig000006ed : STD_LOGIC; 
  signal blk00000003_sig000006ec : STD_LOGIC; 
  signal blk00000003_sig000006eb : STD_LOGIC; 
  signal blk00000003_sig000006ea : STD_LOGIC; 
  signal blk00000003_sig000006e9 : STD_LOGIC; 
  signal blk00000003_sig000006e8 : STD_LOGIC; 
  signal blk00000003_sig000006e7 : STD_LOGIC; 
  signal blk00000003_sig000006e6 : STD_LOGIC; 
  signal blk00000003_sig000006e5 : STD_LOGIC; 
  signal blk00000003_sig000006e4 : STD_LOGIC; 
  signal blk00000003_sig000006e3 : STD_LOGIC; 
  signal blk00000003_sig000006e2 : STD_LOGIC; 
  signal blk00000003_sig000006e1 : STD_LOGIC; 
  signal blk00000003_sig000006e0 : STD_LOGIC; 
  signal blk00000003_sig000006df : STD_LOGIC; 
  signal blk00000003_sig000006de : STD_LOGIC; 
  signal blk00000003_sig000006dd : STD_LOGIC; 
  signal blk00000003_sig000006dc : STD_LOGIC; 
  signal blk00000003_sig000006db : STD_LOGIC; 
  signal blk00000003_sig000006da : STD_LOGIC; 
  signal blk00000003_sig000006d9 : STD_LOGIC; 
  signal blk00000003_sig000006d8 : STD_LOGIC; 
  signal blk00000003_sig000006d7 : STD_LOGIC; 
  signal blk00000003_sig000006d6 : STD_LOGIC; 
  signal blk00000003_sig000006d5 : STD_LOGIC; 
  signal blk00000003_sig000006d4 : STD_LOGIC; 
  signal blk00000003_sig000006d3 : STD_LOGIC; 
  signal blk00000003_sig000006d2 : STD_LOGIC; 
  signal blk00000003_sig000006d1 : STD_LOGIC; 
  signal blk00000003_sig000006d0 : STD_LOGIC; 
  signal blk00000003_sig000006cf : STD_LOGIC; 
  signal blk00000003_sig000006ce : STD_LOGIC; 
  signal blk00000003_sig000006cd : STD_LOGIC; 
  signal blk00000003_sig000006cc : STD_LOGIC; 
  signal blk00000003_sig000006cb : STD_LOGIC; 
  signal blk00000003_sig000006ca : STD_LOGIC; 
  signal blk00000003_sig000006c9 : STD_LOGIC; 
  signal blk00000003_sig000006c8 : STD_LOGIC; 
  signal blk00000003_sig000006c7 : STD_LOGIC; 
  signal blk00000003_sig000006c6 : STD_LOGIC; 
  signal blk00000003_sig000006c5 : STD_LOGIC; 
  signal blk00000003_sig000006c4 : STD_LOGIC; 
  signal blk00000003_sig000006c3 : STD_LOGIC; 
  signal blk00000003_sig000006c2 : STD_LOGIC; 
  signal blk00000003_sig000006c1 : STD_LOGIC; 
  signal blk00000003_sig000006c0 : STD_LOGIC; 
  signal blk00000003_sig000006bf : STD_LOGIC; 
  signal blk00000003_sig000006be : STD_LOGIC; 
  signal blk00000003_sig000006bd : STD_LOGIC; 
  signal blk00000003_sig000006bc : STD_LOGIC; 
  signal blk00000003_sig000006bb : STD_LOGIC; 
  signal blk00000003_sig000006ba : STD_LOGIC; 
  signal blk00000003_sig000006b9 : STD_LOGIC; 
  signal blk00000003_sig000006b8 : STD_LOGIC; 
  signal blk00000003_sig000006b7 : STD_LOGIC; 
  signal blk00000003_sig000006b6 : STD_LOGIC; 
  signal blk00000003_sig000006b5 : STD_LOGIC; 
  signal blk00000003_sig000006b4 : STD_LOGIC; 
  signal blk00000003_sig000006b3 : STD_LOGIC; 
  signal blk00000003_sig000006b2 : STD_LOGIC; 
  signal blk00000003_sig000006b1 : STD_LOGIC; 
  signal blk00000003_sig000006b0 : STD_LOGIC; 
  signal blk00000003_sig000006af : STD_LOGIC; 
  signal blk00000003_sig000006ae : STD_LOGIC; 
  signal blk00000003_sig000006ad : STD_LOGIC; 
  signal blk00000003_sig000006ac : STD_LOGIC; 
  signal blk00000003_sig000006ab : STD_LOGIC; 
  signal blk00000003_sig000006aa : STD_LOGIC; 
  signal blk00000003_sig000006a9 : STD_LOGIC; 
  signal blk00000003_sig000006a8 : STD_LOGIC; 
  signal blk00000003_sig000006a7 : STD_LOGIC; 
  signal blk00000003_sig000006a6 : STD_LOGIC; 
  signal blk00000003_sig000006a5 : STD_LOGIC; 
  signal blk00000003_sig000006a4 : STD_LOGIC; 
  signal blk00000003_sig000006a3 : STD_LOGIC; 
  signal blk00000003_sig000006a2 : STD_LOGIC; 
  signal blk00000003_sig000006a1 : STD_LOGIC; 
  signal blk00000003_sig000006a0 : STD_LOGIC; 
  signal blk00000003_sig0000069f : STD_LOGIC; 
  signal blk00000003_sig0000069e : STD_LOGIC; 
  signal blk00000003_sig0000069d : STD_LOGIC; 
  signal blk00000003_sig0000069c : STD_LOGIC; 
  signal blk00000003_sig0000069b : STD_LOGIC; 
  signal blk00000003_sig0000069a : STD_LOGIC; 
  signal blk00000003_sig00000699 : STD_LOGIC; 
  signal blk00000003_sig00000698 : STD_LOGIC; 
  signal blk00000003_sig00000697 : STD_LOGIC; 
  signal blk00000003_sig00000696 : STD_LOGIC; 
  signal blk00000003_sig00000695 : STD_LOGIC; 
  signal blk00000003_sig00000694 : STD_LOGIC; 
  signal blk00000003_sig00000693 : STD_LOGIC; 
  signal blk00000003_sig00000692 : STD_LOGIC; 
  signal blk00000003_sig00000691 : STD_LOGIC; 
  signal blk00000003_sig00000690 : STD_LOGIC; 
  signal blk00000003_sig0000068f : STD_LOGIC; 
  signal blk00000003_sig0000068e : STD_LOGIC; 
  signal blk00000003_sig0000068d : STD_LOGIC; 
  signal blk00000003_sig0000068c : STD_LOGIC; 
  signal blk00000003_sig0000068b : STD_LOGIC; 
  signal blk00000003_sig0000068a : STD_LOGIC; 
  signal blk00000003_sig00000689 : STD_LOGIC; 
  signal blk00000003_sig00000688 : STD_LOGIC; 
  signal blk00000003_sig00000687 : STD_LOGIC; 
  signal blk00000003_sig00000686 : STD_LOGIC; 
  signal blk00000003_sig00000685 : STD_LOGIC; 
  signal blk00000003_sig00000684 : STD_LOGIC; 
  signal blk00000003_sig00000683 : STD_LOGIC; 
  signal blk00000003_sig00000682 : STD_LOGIC; 
  signal blk00000003_sig00000681 : STD_LOGIC; 
  signal blk00000003_sig00000680 : STD_LOGIC; 
  signal blk00000003_sig0000067f : STD_LOGIC; 
  signal blk00000003_sig0000067e : STD_LOGIC; 
  signal blk00000003_sig0000067d : STD_LOGIC; 
  signal blk00000003_sig0000067c : STD_LOGIC; 
  signal blk00000003_sig0000067b : STD_LOGIC; 
  signal blk00000003_sig0000067a : STD_LOGIC; 
  signal blk00000003_sig00000679 : STD_LOGIC; 
  signal blk00000003_sig00000678 : STD_LOGIC; 
  signal blk00000003_sig00000677 : STD_LOGIC; 
  signal blk00000003_sig00000676 : STD_LOGIC; 
  signal blk00000003_sig00000675 : STD_LOGIC; 
  signal blk00000003_sig00000674 : STD_LOGIC; 
  signal blk00000003_sig00000673 : STD_LOGIC; 
  signal blk00000003_sig00000672 : STD_LOGIC; 
  signal blk00000003_sig00000671 : STD_LOGIC; 
  signal blk00000003_sig00000670 : STD_LOGIC; 
  signal blk00000003_sig0000066f : STD_LOGIC; 
  signal blk00000003_sig0000066e : STD_LOGIC; 
  signal blk00000003_sig0000066d : STD_LOGIC; 
  signal blk00000003_sig0000066c : STD_LOGIC; 
  signal blk00000003_sig0000066b : STD_LOGIC; 
  signal blk00000003_sig0000066a : STD_LOGIC; 
  signal blk00000003_sig00000669 : STD_LOGIC; 
  signal blk00000003_sig00000668 : STD_LOGIC; 
  signal blk00000003_sig00000667 : STD_LOGIC; 
  signal blk00000003_sig00000666 : STD_LOGIC; 
  signal blk00000003_sig00000665 : STD_LOGIC; 
  signal blk00000003_sig00000664 : STD_LOGIC; 
  signal blk00000003_sig00000663 : STD_LOGIC; 
  signal blk00000003_sig00000662 : STD_LOGIC; 
  signal blk00000003_sig00000661 : STD_LOGIC; 
  signal blk00000003_sig00000660 : STD_LOGIC; 
  signal blk00000003_sig0000065f : STD_LOGIC; 
  signal blk00000003_sig0000065e : STD_LOGIC; 
  signal blk00000003_sig0000065d : STD_LOGIC; 
  signal blk00000003_sig0000065c : STD_LOGIC; 
  signal blk00000003_sig0000065b : STD_LOGIC; 
  signal blk00000003_sig0000065a : STD_LOGIC; 
  signal blk00000003_sig00000659 : STD_LOGIC; 
  signal blk00000003_sig00000658 : STD_LOGIC; 
  signal blk00000003_sig00000657 : STD_LOGIC; 
  signal blk00000003_sig00000656 : STD_LOGIC; 
  signal blk00000003_sig00000655 : STD_LOGIC; 
  signal blk00000003_sig00000654 : STD_LOGIC; 
  signal blk00000003_sig00000653 : STD_LOGIC; 
  signal blk00000003_sig00000652 : STD_LOGIC; 
  signal blk00000003_sig00000651 : STD_LOGIC; 
  signal blk00000003_sig00000650 : STD_LOGIC; 
  signal blk00000003_sig0000064f : STD_LOGIC; 
  signal blk00000003_sig0000064e : STD_LOGIC; 
  signal blk00000003_sig0000064d : STD_LOGIC; 
  signal blk00000003_sig0000064c : STD_LOGIC; 
  signal blk00000003_sig0000064b : STD_LOGIC; 
  signal blk00000003_sig0000064a : STD_LOGIC; 
  signal blk00000003_sig00000649 : STD_LOGIC; 
  signal blk00000003_sig00000648 : STD_LOGIC; 
  signal blk00000003_sig00000647 : STD_LOGIC; 
  signal blk00000003_sig00000646 : STD_LOGIC; 
  signal blk00000003_sig00000645 : STD_LOGIC; 
  signal blk00000003_sig00000644 : STD_LOGIC; 
  signal blk00000003_sig00000643 : STD_LOGIC; 
  signal blk00000003_sig00000642 : STD_LOGIC; 
  signal blk00000003_sig00000641 : STD_LOGIC; 
  signal blk00000003_sig00000640 : STD_LOGIC; 
  signal blk00000003_sig0000063f : STD_LOGIC; 
  signal blk00000003_sig0000063e : STD_LOGIC; 
  signal blk00000003_sig0000063d : STD_LOGIC; 
  signal blk00000003_sig0000063c : STD_LOGIC; 
  signal blk00000003_sig0000063b : STD_LOGIC; 
  signal blk00000003_sig0000063a : STD_LOGIC; 
  signal blk00000003_sig00000639 : STD_LOGIC; 
  signal blk00000003_sig00000638 : STD_LOGIC; 
  signal blk00000003_sig00000637 : STD_LOGIC; 
  signal blk00000003_sig00000636 : STD_LOGIC; 
  signal blk00000003_sig00000635 : STD_LOGIC; 
  signal blk00000003_sig00000634 : STD_LOGIC; 
  signal blk00000003_sig00000633 : STD_LOGIC; 
  signal blk00000003_sig00000632 : STD_LOGIC; 
  signal blk00000003_sig00000631 : STD_LOGIC; 
  signal blk00000003_sig00000630 : STD_LOGIC; 
  signal blk00000003_sig0000062f : STD_LOGIC; 
  signal blk00000003_sig0000062e : STD_LOGIC; 
  signal blk00000003_sig0000062d : STD_LOGIC; 
  signal blk00000003_sig0000062c : STD_LOGIC; 
  signal blk00000003_sig0000062b : STD_LOGIC; 
  signal blk00000003_sig0000062a : STD_LOGIC; 
  signal blk00000003_sig00000629 : STD_LOGIC; 
  signal blk00000003_sig00000628 : STD_LOGIC; 
  signal blk00000003_sig00000627 : STD_LOGIC; 
  signal blk00000003_sig00000626 : STD_LOGIC; 
  signal blk00000003_sig00000625 : STD_LOGIC; 
  signal blk00000003_sig00000624 : STD_LOGIC; 
  signal blk00000003_sig00000623 : STD_LOGIC; 
  signal blk00000003_sig00000622 : STD_LOGIC; 
  signal blk00000003_sig00000621 : STD_LOGIC; 
  signal blk00000003_sig00000620 : STD_LOGIC; 
  signal blk00000003_sig0000061f : STD_LOGIC; 
  signal blk00000003_sig0000061e : STD_LOGIC; 
  signal blk00000003_sig0000061d : STD_LOGIC; 
  signal blk00000003_sig0000061c : STD_LOGIC; 
  signal blk00000003_sig0000061b : STD_LOGIC; 
  signal blk00000003_sig0000061a : STD_LOGIC; 
  signal blk00000003_sig00000619 : STD_LOGIC; 
  signal blk00000003_sig00000618 : STD_LOGIC; 
  signal blk00000003_sig00000617 : STD_LOGIC; 
  signal blk00000003_sig00000616 : STD_LOGIC; 
  signal blk00000003_sig00000615 : STD_LOGIC; 
  signal blk00000003_sig00000614 : STD_LOGIC; 
  signal blk00000003_sig00000613 : STD_LOGIC; 
  signal blk00000003_sig00000612 : STD_LOGIC; 
  signal blk00000003_sig00000611 : STD_LOGIC; 
  signal blk00000003_sig00000610 : STD_LOGIC; 
  signal blk00000003_sig0000060f : STD_LOGIC; 
  signal blk00000003_sig0000060e : STD_LOGIC; 
  signal blk00000003_sig0000060d : STD_LOGIC; 
  signal blk00000003_sig0000060c : STD_LOGIC; 
  signal blk00000003_sig0000060b : STD_LOGIC; 
  signal blk00000003_sig0000060a : STD_LOGIC; 
  signal blk00000003_sig00000609 : STD_LOGIC; 
  signal blk00000003_sig00000608 : STD_LOGIC; 
  signal blk00000003_sig00000607 : STD_LOGIC; 
  signal blk00000003_sig00000606 : STD_LOGIC; 
  signal blk00000003_sig00000605 : STD_LOGIC; 
  signal blk00000003_sig00000604 : STD_LOGIC; 
  signal blk00000003_sig00000603 : STD_LOGIC; 
  signal blk00000003_sig00000602 : STD_LOGIC; 
  signal blk00000003_sig00000601 : STD_LOGIC; 
  signal blk00000003_sig00000600 : STD_LOGIC; 
  signal blk00000003_sig000005ff : STD_LOGIC; 
  signal blk00000003_sig000005fe : STD_LOGIC; 
  signal blk00000003_sig000005fd : STD_LOGIC; 
  signal blk00000003_sig000005fc : STD_LOGIC; 
  signal blk00000003_sig000005fb : STD_LOGIC; 
  signal blk00000003_sig000005fa : STD_LOGIC; 
  signal blk00000003_sig000005f9 : STD_LOGIC; 
  signal blk00000003_sig000005f8 : STD_LOGIC; 
  signal blk00000003_sig000005f7 : STD_LOGIC; 
  signal blk00000003_sig000005f6 : STD_LOGIC; 
  signal blk00000003_sig000005f5 : STD_LOGIC; 
  signal blk00000003_sig000005f4 : STD_LOGIC; 
  signal blk00000003_sig000005f3 : STD_LOGIC; 
  signal blk00000003_sig000005f2 : STD_LOGIC; 
  signal blk00000003_sig000005f1 : STD_LOGIC; 
  signal blk00000003_sig000005f0 : STD_LOGIC; 
  signal blk00000003_sig000005ef : STD_LOGIC; 
  signal blk00000003_sig000005ee : STD_LOGIC; 
  signal blk00000003_sig000005ed : STD_LOGIC; 
  signal blk00000003_sig000005ec : STD_LOGIC; 
  signal blk00000003_sig000005eb : STD_LOGIC; 
  signal blk00000003_sig000005ea : STD_LOGIC; 
  signal blk00000003_sig000005e9 : STD_LOGIC; 
  signal blk00000003_sig000005e8 : STD_LOGIC; 
  signal blk00000003_sig000005e7 : STD_LOGIC; 
  signal blk00000003_sig000005e6 : STD_LOGIC; 
  signal blk00000003_sig000005e5 : STD_LOGIC; 
  signal blk00000003_sig000005e4 : STD_LOGIC; 
  signal blk00000003_sig000005e3 : STD_LOGIC; 
  signal blk00000003_sig000005e2 : STD_LOGIC; 
  signal blk00000003_sig000005e1 : STD_LOGIC; 
  signal blk00000003_sig000005e0 : STD_LOGIC; 
  signal blk00000003_sig000005df : STD_LOGIC; 
  signal blk00000003_sig000005de : STD_LOGIC; 
  signal blk00000003_sig000005dd : STD_LOGIC; 
  signal blk00000003_sig000005dc : STD_LOGIC; 
  signal blk00000003_sig000005db : STD_LOGIC; 
  signal blk00000003_sig000005da : STD_LOGIC; 
  signal blk00000003_sig000005d9 : STD_LOGIC; 
  signal blk00000003_sig000005d8 : STD_LOGIC; 
  signal blk00000003_sig000005d7 : STD_LOGIC; 
  signal blk00000003_sig000005d6 : STD_LOGIC; 
  signal blk00000003_sig000005d5 : STD_LOGIC; 
  signal blk00000003_sig000005d4 : STD_LOGIC; 
  signal blk00000003_sig000005d3 : STD_LOGIC; 
  signal blk00000003_sig000005d2 : STD_LOGIC; 
  signal blk00000003_sig000005d1 : STD_LOGIC; 
  signal blk00000003_sig000005d0 : STD_LOGIC; 
  signal blk00000003_sig000005cf : STD_LOGIC; 
  signal blk00000003_sig000005ce : STD_LOGIC; 
  signal blk00000003_sig000005cd : STD_LOGIC; 
  signal blk00000003_sig000005cc : STD_LOGIC; 
  signal blk00000003_sig000005cb : STD_LOGIC; 
  signal blk00000003_sig000005ca : STD_LOGIC; 
  signal blk00000003_sig000005c9 : STD_LOGIC; 
  signal blk00000003_sig000005c8 : STD_LOGIC; 
  signal blk00000003_sig000005c7 : STD_LOGIC; 
  signal blk00000003_sig000005c6 : STD_LOGIC; 
  signal blk00000003_sig000005c5 : STD_LOGIC; 
  signal blk00000003_sig000005c4 : STD_LOGIC; 
  signal blk00000003_sig000005c3 : STD_LOGIC; 
  signal blk00000003_sig000005c2 : STD_LOGIC; 
  signal blk00000003_sig000005c1 : STD_LOGIC; 
  signal blk00000003_sig000005c0 : STD_LOGIC; 
  signal blk00000003_sig000005bf : STD_LOGIC; 
  signal blk00000003_sig000005be : STD_LOGIC; 
  signal blk00000003_sig000005bd : STD_LOGIC; 
  signal blk00000003_sig000005bc : STD_LOGIC; 
  signal blk00000003_sig000005bb : STD_LOGIC; 
  signal blk00000003_sig000005ba : STD_LOGIC; 
  signal blk00000003_sig000005b9 : STD_LOGIC; 
  signal blk00000003_sig000005b8 : STD_LOGIC; 
  signal blk00000003_sig000005b7 : STD_LOGIC; 
  signal blk00000003_sig000005b6 : STD_LOGIC; 
  signal blk00000003_sig000005b5 : STD_LOGIC; 
  signal blk00000003_sig000005b4 : STD_LOGIC; 
  signal blk00000003_sig000005b3 : STD_LOGIC; 
  signal blk00000003_sig000005b2 : STD_LOGIC; 
  signal blk00000003_sig000005b1 : STD_LOGIC; 
  signal blk00000003_sig000005b0 : STD_LOGIC; 
  signal blk00000003_sig000005af : STD_LOGIC; 
  signal blk00000003_sig000005ae : STD_LOGIC; 
  signal blk00000003_sig000005ad : STD_LOGIC; 
  signal blk00000003_sig000005ac : STD_LOGIC; 
  signal blk00000003_sig000005ab : STD_LOGIC; 
  signal blk00000003_sig000005aa : STD_LOGIC; 
  signal blk00000003_sig000005a9 : STD_LOGIC; 
  signal blk00000003_sig000005a8 : STD_LOGIC; 
  signal blk00000003_sig000005a7 : STD_LOGIC; 
  signal blk00000003_sig000005a6 : STD_LOGIC; 
  signal blk00000003_sig000005a5 : STD_LOGIC; 
  signal blk00000003_sig000005a4 : STD_LOGIC; 
  signal blk00000003_sig000005a3 : STD_LOGIC; 
  signal blk00000003_sig000005a2 : STD_LOGIC; 
  signal blk00000003_sig000005a1 : STD_LOGIC; 
  signal blk00000003_sig000005a0 : STD_LOGIC; 
  signal blk00000003_sig0000059f : STD_LOGIC; 
  signal blk00000003_sig0000059e : STD_LOGIC; 
  signal blk00000003_sig0000059d : STD_LOGIC; 
  signal blk00000003_sig0000059c : STD_LOGIC; 
  signal blk00000003_sig0000059b : STD_LOGIC; 
  signal blk00000003_sig0000059a : STD_LOGIC; 
  signal blk00000003_sig00000599 : STD_LOGIC; 
  signal blk00000003_sig00000598 : STD_LOGIC; 
  signal blk00000003_sig00000597 : STD_LOGIC; 
  signal blk00000003_sig00000596 : STD_LOGIC; 
  signal blk00000003_sig00000595 : STD_LOGIC; 
  signal blk00000003_sig00000594 : STD_LOGIC; 
  signal blk00000003_sig00000593 : STD_LOGIC; 
  signal blk00000003_sig00000592 : STD_LOGIC; 
  signal blk00000003_sig00000591 : STD_LOGIC; 
  signal blk00000003_sig00000590 : STD_LOGIC; 
  signal blk00000003_sig0000058f : STD_LOGIC; 
  signal blk00000003_sig0000058e : STD_LOGIC; 
  signal blk00000003_sig0000058d : STD_LOGIC; 
  signal blk00000003_sig0000058c : STD_LOGIC; 
  signal blk00000003_sig0000058b : STD_LOGIC; 
  signal blk00000003_sig0000058a : STD_LOGIC; 
  signal blk00000003_sig00000589 : STD_LOGIC; 
  signal blk00000003_sig00000588 : STD_LOGIC; 
  signal blk00000003_sig00000587 : STD_LOGIC; 
  signal blk00000003_sig00000586 : STD_LOGIC; 
  signal blk00000003_sig00000585 : STD_LOGIC; 
  signal blk00000003_sig00000584 : STD_LOGIC; 
  signal blk00000003_sig00000583 : STD_LOGIC; 
  signal blk00000003_sig00000582 : STD_LOGIC; 
  signal blk00000003_sig00000581 : STD_LOGIC; 
  signal blk00000003_sig00000580 : STD_LOGIC; 
  signal blk00000003_sig0000057f : STD_LOGIC; 
  signal blk00000003_sig0000057e : STD_LOGIC; 
  signal blk00000003_sig0000057d : STD_LOGIC; 
  signal blk00000003_sig0000057c : STD_LOGIC; 
  signal blk00000003_sig0000057b : STD_LOGIC; 
  signal blk00000003_sig0000057a : STD_LOGIC; 
  signal blk00000003_sig00000579 : STD_LOGIC; 
  signal blk00000003_sig00000578 : STD_LOGIC; 
  signal blk00000003_sig00000577 : STD_LOGIC; 
  signal blk00000003_sig00000576 : STD_LOGIC; 
  signal blk00000003_sig00000575 : STD_LOGIC; 
  signal blk00000003_sig00000574 : STD_LOGIC; 
  signal blk00000003_sig00000573 : STD_LOGIC; 
  signal blk00000003_sig00000572 : STD_LOGIC; 
  signal blk00000003_sig00000571 : STD_LOGIC; 
  signal blk00000003_sig00000570 : STD_LOGIC; 
  signal blk00000003_sig0000056f : STD_LOGIC; 
  signal blk00000003_sig0000056e : STD_LOGIC; 
  signal blk00000003_sig0000056d : STD_LOGIC; 
  signal blk00000003_sig0000056c : STD_LOGIC; 
  signal blk00000003_sig0000056b : STD_LOGIC; 
  signal blk00000003_sig0000056a : STD_LOGIC; 
  signal blk00000003_sig00000569 : STD_LOGIC; 
  signal blk00000003_sig00000568 : STD_LOGIC; 
  signal blk00000003_sig00000567 : STD_LOGIC; 
  signal blk00000003_sig00000566 : STD_LOGIC; 
  signal blk00000003_sig00000565 : STD_LOGIC; 
  signal blk00000003_sig00000564 : STD_LOGIC; 
  signal blk00000003_sig00000563 : STD_LOGIC; 
  signal blk00000003_sig00000562 : STD_LOGIC; 
  signal blk00000003_sig00000561 : STD_LOGIC; 
  signal blk00000003_sig00000560 : STD_LOGIC; 
  signal blk00000003_sig0000055f : STD_LOGIC; 
  signal blk00000003_sig0000055e : STD_LOGIC; 
  signal blk00000003_sig0000055d : STD_LOGIC; 
  signal blk00000003_sig0000055c : STD_LOGIC; 
  signal blk00000003_sig0000055b : STD_LOGIC; 
  signal blk00000003_sig0000055a : STD_LOGIC; 
  signal blk00000003_sig00000559 : STD_LOGIC; 
  signal blk00000003_sig00000558 : STD_LOGIC; 
  signal blk00000003_sig00000557 : STD_LOGIC; 
  signal blk00000003_sig00000556 : STD_LOGIC; 
  signal blk00000003_sig00000555 : STD_LOGIC; 
  signal blk00000003_sig00000554 : STD_LOGIC; 
  signal blk00000003_sig00000553 : STD_LOGIC; 
  signal blk00000003_sig00000552 : STD_LOGIC; 
  signal blk00000003_sig00000551 : STD_LOGIC; 
  signal blk00000003_sig00000550 : STD_LOGIC; 
  signal blk00000003_sig0000054f : STD_LOGIC; 
  signal blk00000003_sig0000054e : STD_LOGIC; 
  signal blk00000003_sig0000054d : STD_LOGIC; 
  signal blk00000003_sig0000054c : STD_LOGIC; 
  signal blk00000003_sig0000054b : STD_LOGIC; 
  signal blk00000003_sig0000054a : STD_LOGIC; 
  signal blk00000003_sig00000549 : STD_LOGIC; 
  signal blk00000003_sig00000548 : STD_LOGIC; 
  signal blk00000003_sig00000547 : STD_LOGIC; 
  signal blk00000003_sig00000546 : STD_LOGIC; 
  signal blk00000003_sig00000545 : STD_LOGIC; 
  signal blk00000003_sig00000544 : STD_LOGIC; 
  signal blk00000003_sig00000543 : STD_LOGIC; 
  signal blk00000003_sig00000542 : STD_LOGIC; 
  signal blk00000003_sig00000541 : STD_LOGIC; 
  signal blk00000003_sig00000540 : STD_LOGIC; 
  signal blk00000003_sig0000053f : STD_LOGIC; 
  signal blk00000003_sig0000053e : STD_LOGIC; 
  signal blk00000003_sig0000053d : STD_LOGIC; 
  signal blk00000003_sig0000053c : STD_LOGIC; 
  signal blk00000003_sig0000053b : STD_LOGIC; 
  signal blk00000003_sig0000053a : STD_LOGIC; 
  signal blk00000003_sig00000539 : STD_LOGIC; 
  signal blk00000003_sig00000538 : STD_LOGIC; 
  signal blk00000003_sig00000537 : STD_LOGIC; 
  signal blk00000003_sig00000536 : STD_LOGIC; 
  signal blk00000003_sig00000535 : STD_LOGIC; 
  signal blk00000003_sig00000534 : STD_LOGIC; 
  signal blk00000003_sig00000533 : STD_LOGIC; 
  signal blk00000003_sig00000532 : STD_LOGIC; 
  signal blk00000003_sig00000531 : STD_LOGIC; 
  signal blk00000003_sig00000530 : STD_LOGIC; 
  signal blk00000003_sig0000052f : STD_LOGIC; 
  signal blk00000003_sig0000052e : STD_LOGIC; 
  signal blk00000003_sig0000052d : STD_LOGIC; 
  signal blk00000003_sig0000052c : STD_LOGIC; 
  signal blk00000003_sig0000052b : STD_LOGIC; 
  signal blk00000003_sig0000052a : STD_LOGIC; 
  signal blk00000003_sig00000529 : STD_LOGIC; 
  signal blk00000003_sig00000528 : STD_LOGIC; 
  signal blk00000003_sig00000527 : STD_LOGIC; 
  signal blk00000003_sig00000526 : STD_LOGIC; 
  signal blk00000003_sig00000525 : STD_LOGIC; 
  signal blk00000003_sig00000524 : STD_LOGIC; 
  signal blk00000003_sig00000523 : STD_LOGIC; 
  signal blk00000003_sig00000522 : STD_LOGIC; 
  signal blk00000003_sig00000521 : STD_LOGIC; 
  signal blk00000003_sig00000520 : STD_LOGIC; 
  signal blk00000003_sig0000051f : STD_LOGIC; 
  signal blk00000003_sig0000051e : STD_LOGIC; 
  signal blk00000003_sig0000051d : STD_LOGIC; 
  signal blk00000003_sig0000051c : STD_LOGIC; 
  signal blk00000003_sig0000051b : STD_LOGIC; 
  signal blk00000003_sig0000051a : STD_LOGIC; 
  signal blk00000003_sig00000519 : STD_LOGIC; 
  signal blk00000003_sig00000518 : STD_LOGIC; 
  signal blk00000003_sig00000517 : STD_LOGIC; 
  signal blk00000003_sig00000516 : STD_LOGIC; 
  signal blk00000003_sig00000515 : STD_LOGIC; 
  signal blk00000003_sig00000514 : STD_LOGIC; 
  signal blk00000003_sig00000513 : STD_LOGIC; 
  signal blk00000003_sig00000512 : STD_LOGIC; 
  signal blk00000003_sig00000511 : STD_LOGIC; 
  signal blk00000003_sig00000510 : STD_LOGIC; 
  signal blk00000003_sig0000050f : STD_LOGIC; 
  signal blk00000003_sig0000050e : STD_LOGIC; 
  signal blk00000003_sig0000050d : STD_LOGIC; 
  signal blk00000003_sig0000050c : STD_LOGIC; 
  signal blk00000003_sig0000050b : STD_LOGIC; 
  signal blk00000003_sig0000050a : STD_LOGIC; 
  signal blk00000003_sig00000509 : STD_LOGIC; 
  signal blk00000003_sig00000508 : STD_LOGIC; 
  signal blk00000003_sig00000507 : STD_LOGIC; 
  signal blk00000003_sig00000506 : STD_LOGIC; 
  signal blk00000003_sig00000505 : STD_LOGIC; 
  signal blk00000003_sig00000504 : STD_LOGIC; 
  signal blk00000003_sig00000503 : STD_LOGIC; 
  signal blk00000003_sig00000502 : STD_LOGIC; 
  signal blk00000003_sig00000501 : STD_LOGIC; 
  signal blk00000003_sig00000500 : STD_LOGIC; 
  signal blk00000003_sig000004ff : STD_LOGIC; 
  signal blk00000003_sig000004fe : STD_LOGIC; 
  signal blk00000003_sig000004fd : STD_LOGIC; 
  signal blk00000003_sig000004fc : STD_LOGIC; 
  signal blk00000003_sig000004fb : STD_LOGIC; 
  signal blk00000003_sig000004fa : STD_LOGIC; 
  signal blk00000003_sig000004f9 : STD_LOGIC; 
  signal blk00000003_sig000004f8 : STD_LOGIC; 
  signal blk00000003_sig000004f7 : STD_LOGIC; 
  signal blk00000003_sig000004f6 : STD_LOGIC; 
  signal blk00000003_sig000004f5 : STD_LOGIC; 
  signal blk00000003_sig000004f4 : STD_LOGIC; 
  signal blk00000003_sig000004f3 : STD_LOGIC; 
  signal blk00000003_sig000004f2 : STD_LOGIC; 
  signal blk00000003_sig000004f1 : STD_LOGIC; 
  signal blk00000003_sig000004f0 : STD_LOGIC; 
  signal blk00000003_sig000004ef : STD_LOGIC; 
  signal blk00000003_sig000004ee : STD_LOGIC; 
  signal blk00000003_sig000004ed : STD_LOGIC; 
  signal blk00000003_sig000004ec : STD_LOGIC; 
  signal blk00000003_sig000004eb : STD_LOGIC; 
  signal blk00000003_sig000004ea : STD_LOGIC; 
  signal blk00000003_sig000004e9 : STD_LOGIC; 
  signal blk00000003_sig000004e8 : STD_LOGIC; 
  signal blk00000003_sig000004e7 : STD_LOGIC; 
  signal blk00000003_sig000004e6 : STD_LOGIC; 
  signal blk00000003_sig000004e5 : STD_LOGIC; 
  signal blk00000003_sig000004e4 : STD_LOGIC; 
  signal blk00000003_sig000004e3 : STD_LOGIC; 
  signal blk00000003_sig000004e2 : STD_LOGIC; 
  signal blk00000003_sig000004e1 : STD_LOGIC; 
  signal blk00000003_sig000004e0 : STD_LOGIC; 
  signal blk00000003_sig000004df : STD_LOGIC; 
  signal blk00000003_sig000004de : STD_LOGIC; 
  signal blk00000003_sig000004dd : STD_LOGIC; 
  signal blk00000003_sig000004dc : STD_LOGIC; 
  signal blk00000003_sig000004db : STD_LOGIC; 
  signal blk00000003_sig000004da : STD_LOGIC; 
  signal blk00000003_sig000004d9 : STD_LOGIC; 
  signal blk00000003_sig000004d8 : STD_LOGIC; 
  signal blk00000003_sig000004d7 : STD_LOGIC; 
  signal blk00000003_sig000004d6 : STD_LOGIC; 
  signal blk00000003_sig000004d5 : STD_LOGIC; 
  signal blk00000003_sig000004d4 : STD_LOGIC; 
  signal blk00000003_sig000004d3 : STD_LOGIC; 
  signal blk00000003_sig000004d2 : STD_LOGIC; 
  signal blk00000003_sig000004d1 : STD_LOGIC; 
  signal blk00000003_sig000004d0 : STD_LOGIC; 
  signal blk00000003_sig000004cf : STD_LOGIC; 
  signal blk00000003_sig000004ce : STD_LOGIC; 
  signal blk00000003_sig000004cd : STD_LOGIC; 
  signal blk00000003_sig000004cc : STD_LOGIC; 
  signal blk00000003_sig000004cb : STD_LOGIC; 
  signal blk00000003_sig000004ca : STD_LOGIC; 
  signal blk00000003_sig000004c9 : STD_LOGIC; 
  signal blk00000003_sig000004c8 : STD_LOGIC; 
  signal blk00000003_sig000004c7 : STD_LOGIC; 
  signal blk00000003_sig000004c6 : STD_LOGIC; 
  signal blk00000003_sig000004c5 : STD_LOGIC; 
  signal blk00000003_sig000004c4 : STD_LOGIC; 
  signal blk00000003_sig000004c3 : STD_LOGIC; 
  signal blk00000003_sig000004c2 : STD_LOGIC; 
  signal blk00000003_sig000004c1 : STD_LOGIC; 
  signal blk00000003_sig000004c0 : STD_LOGIC; 
  signal blk00000003_sig000004bf : STD_LOGIC; 
  signal blk00000003_sig000004be : STD_LOGIC; 
  signal blk00000003_sig000004bd : STD_LOGIC; 
  signal blk00000003_sig000004bc : STD_LOGIC; 
  signal blk00000003_sig000004bb : STD_LOGIC; 
  signal blk00000003_sig000004ba : STD_LOGIC; 
  signal blk00000003_sig000004b9 : STD_LOGIC; 
  signal blk00000003_sig000004b8 : STD_LOGIC; 
  signal blk00000003_sig000004b7 : STD_LOGIC; 
  signal blk00000003_sig000004b6 : STD_LOGIC; 
  signal blk00000003_sig000004b5 : STD_LOGIC; 
  signal blk00000003_sig000004b4 : STD_LOGIC; 
  signal blk00000003_sig000004b3 : STD_LOGIC; 
  signal blk00000003_sig000004b2 : STD_LOGIC; 
  signal blk00000003_sig000004b1 : STD_LOGIC; 
  signal blk00000003_sig000004b0 : STD_LOGIC; 
  signal blk00000003_sig000004af : STD_LOGIC; 
  signal blk00000003_sig000004ae : STD_LOGIC; 
  signal blk00000003_sig000004ad : STD_LOGIC; 
  signal blk00000003_sig000004ac : STD_LOGIC; 
  signal blk00000003_sig000004ab : STD_LOGIC; 
  signal blk00000003_sig000004aa : STD_LOGIC; 
  signal blk00000003_sig000004a9 : STD_LOGIC; 
  signal blk00000003_sig000004a8 : STD_LOGIC; 
  signal blk00000003_sig000004a7 : STD_LOGIC; 
  signal blk00000003_sig000004a6 : STD_LOGIC; 
  signal blk00000003_sig000004a5 : STD_LOGIC; 
  signal blk00000003_sig000004a4 : STD_LOGIC; 
  signal blk00000003_sig000004a3 : STD_LOGIC; 
  signal blk00000003_sig000004a2 : STD_LOGIC; 
  signal blk00000003_sig000004a1 : STD_LOGIC; 
  signal blk00000003_sig000004a0 : STD_LOGIC; 
  signal blk00000003_sig0000049f : STD_LOGIC; 
  signal blk00000003_sig0000049e : STD_LOGIC; 
  signal blk00000003_sig0000049d : STD_LOGIC; 
  signal blk00000003_sig0000049c : STD_LOGIC; 
  signal blk00000003_sig0000049b : STD_LOGIC; 
  signal blk00000003_sig0000049a : STD_LOGIC; 
  signal blk00000003_sig00000499 : STD_LOGIC; 
  signal blk00000003_sig00000498 : STD_LOGIC; 
  signal blk00000003_sig00000497 : STD_LOGIC; 
  signal blk00000003_sig00000496 : STD_LOGIC; 
  signal blk00000003_sig00000495 : STD_LOGIC; 
  signal blk00000003_sig00000494 : STD_LOGIC; 
  signal blk00000003_sig00000493 : STD_LOGIC; 
  signal blk00000003_sig00000492 : STD_LOGIC; 
  signal blk00000003_sig00000491 : STD_LOGIC; 
  signal blk00000003_sig00000490 : STD_LOGIC; 
  signal blk00000003_sig0000048f : STD_LOGIC; 
  signal blk00000003_sig0000048e : STD_LOGIC; 
  signal blk00000003_sig0000048d : STD_LOGIC; 
  signal blk00000003_sig0000048c : STD_LOGIC; 
  signal blk00000003_sig0000048b : STD_LOGIC; 
  signal blk00000003_sig0000048a : STD_LOGIC; 
  signal blk00000003_sig00000489 : STD_LOGIC; 
  signal blk00000003_sig00000488 : STD_LOGIC; 
  signal blk00000003_sig00000487 : STD_LOGIC; 
  signal blk00000003_sig00000486 : STD_LOGIC; 
  signal blk00000003_sig00000485 : STD_LOGIC; 
  signal blk00000003_sig00000484 : STD_LOGIC; 
  signal blk00000003_sig00000483 : STD_LOGIC; 
  signal blk00000003_sig00000482 : STD_LOGIC; 
  signal blk00000003_sig00000481 : STD_LOGIC; 
  signal blk00000003_sig00000480 : STD_LOGIC; 
  signal blk00000003_sig0000047f : STD_LOGIC; 
  signal blk00000003_sig0000047e : STD_LOGIC; 
  signal blk00000003_sig0000047d : STD_LOGIC; 
  signal blk00000003_sig0000047c : STD_LOGIC; 
  signal blk00000003_sig0000047b : STD_LOGIC; 
  signal blk00000003_sig0000047a : STD_LOGIC; 
  signal blk00000003_sig00000479 : STD_LOGIC; 
  signal blk00000003_sig00000478 : STD_LOGIC; 
  signal blk00000003_sig00000477 : STD_LOGIC; 
  signal blk00000003_sig00000476 : STD_LOGIC; 
  signal blk00000003_sig00000475 : STD_LOGIC; 
  signal blk00000003_sig00000474 : STD_LOGIC; 
  signal blk00000003_sig00000473 : STD_LOGIC; 
  signal blk00000003_sig00000472 : STD_LOGIC; 
  signal blk00000003_sig00000471 : STD_LOGIC; 
  signal blk00000003_sig00000470 : STD_LOGIC; 
  signal blk00000003_sig0000046f : STD_LOGIC; 
  signal blk00000003_sig0000046e : STD_LOGIC; 
  signal blk00000003_sig0000046d : STD_LOGIC; 
  signal blk00000003_sig0000046c : STD_LOGIC; 
  signal blk00000003_sig0000046b : STD_LOGIC; 
  signal blk00000003_sig0000046a : STD_LOGIC; 
  signal blk00000003_sig00000469 : STD_LOGIC; 
  signal blk00000003_sig00000468 : STD_LOGIC; 
  signal blk00000003_sig00000467 : STD_LOGIC; 
  signal blk00000003_sig00000466 : STD_LOGIC; 
  signal blk00000003_sig00000465 : STD_LOGIC; 
  signal blk00000003_sig00000464 : STD_LOGIC; 
  signal blk00000003_sig00000463 : STD_LOGIC; 
  signal blk00000003_sig00000462 : STD_LOGIC; 
  signal blk00000003_sig00000461 : STD_LOGIC; 
  signal blk00000003_sig00000460 : STD_LOGIC; 
  signal blk00000003_sig0000045f : STD_LOGIC; 
  signal blk00000003_sig0000045e : STD_LOGIC; 
  signal blk00000003_sig0000045d : STD_LOGIC; 
  signal blk00000003_sig0000045c : STD_LOGIC; 
  signal blk00000003_sig0000045b : STD_LOGIC; 
  signal blk00000003_sig0000045a : STD_LOGIC; 
  signal blk00000003_sig00000459 : STD_LOGIC; 
  signal blk00000003_sig00000458 : STD_LOGIC; 
  signal blk00000003_sig00000457 : STD_LOGIC; 
  signal blk00000003_sig00000456 : STD_LOGIC; 
  signal blk00000003_sig00000455 : STD_LOGIC; 
  signal blk00000003_sig00000454 : STD_LOGIC; 
  signal blk00000003_sig00000453 : STD_LOGIC; 
  signal blk00000003_sig00000452 : STD_LOGIC; 
  signal blk00000003_sig00000451 : STD_LOGIC; 
  signal blk00000003_sig00000450 : STD_LOGIC; 
  signal blk00000003_sig0000044f : STD_LOGIC; 
  signal blk00000003_sig0000044e : STD_LOGIC; 
  signal blk00000003_sig0000044d : STD_LOGIC; 
  signal blk00000003_sig0000044c : STD_LOGIC; 
  signal blk00000003_sig0000044b : STD_LOGIC; 
  signal blk00000003_sig0000044a : STD_LOGIC; 
  signal blk00000003_sig00000449 : STD_LOGIC; 
  signal blk00000003_sig00000448 : STD_LOGIC; 
  signal blk00000003_sig00000447 : STD_LOGIC; 
  signal blk00000003_sig00000446 : STD_LOGIC; 
  signal blk00000003_sig00000445 : STD_LOGIC; 
  signal blk00000003_sig00000444 : STD_LOGIC; 
  signal blk00000003_sig00000443 : STD_LOGIC; 
  signal blk00000003_sig00000442 : STD_LOGIC; 
  signal blk00000003_sig00000441 : STD_LOGIC; 
  signal blk00000003_sig00000440 : STD_LOGIC; 
  signal blk00000003_sig0000043f : STD_LOGIC; 
  signal blk00000003_sig0000043e : STD_LOGIC; 
  signal blk00000003_sig0000043d : STD_LOGIC; 
  signal blk00000003_sig0000043c : STD_LOGIC; 
  signal blk00000003_sig0000043b : STD_LOGIC; 
  signal blk00000003_sig0000043a : STD_LOGIC; 
  signal blk00000003_sig00000439 : STD_LOGIC; 
  signal blk00000003_sig00000438 : STD_LOGIC; 
  signal blk00000003_sig00000437 : STD_LOGIC; 
  signal blk00000003_sig00000436 : STD_LOGIC; 
  signal blk00000003_sig00000435 : STD_LOGIC; 
  signal blk00000003_sig00000434 : STD_LOGIC; 
  signal blk00000003_sig00000433 : STD_LOGIC; 
  signal blk00000003_sig00000432 : STD_LOGIC; 
  signal blk00000003_sig00000431 : STD_LOGIC; 
  signal blk00000003_sig00000430 : STD_LOGIC; 
  signal blk00000003_sig0000042f : STD_LOGIC; 
  signal blk00000003_sig0000042e : STD_LOGIC; 
  signal blk00000003_sig0000042d : STD_LOGIC; 
  signal blk00000003_sig0000042c : STD_LOGIC; 
  signal blk00000003_sig0000042b : STD_LOGIC; 
  signal blk00000003_sig0000042a : STD_LOGIC; 
  signal blk00000003_sig00000429 : STD_LOGIC; 
  signal blk00000003_sig00000428 : STD_LOGIC; 
  signal blk00000003_sig00000427 : STD_LOGIC; 
  signal blk00000003_sig00000426 : STD_LOGIC; 
  signal blk00000003_sig00000425 : STD_LOGIC; 
  signal blk00000003_sig00000424 : STD_LOGIC; 
  signal blk00000003_sig00000423 : STD_LOGIC; 
  signal blk00000003_sig00000422 : STD_LOGIC; 
  signal blk00000003_sig00000421 : STD_LOGIC; 
  signal blk00000003_sig00000420 : STD_LOGIC; 
  signal blk00000003_sig0000041f : STD_LOGIC; 
  signal blk00000003_sig0000041e : STD_LOGIC; 
  signal blk00000003_sig0000041d : STD_LOGIC; 
  signal blk00000003_sig0000041c : STD_LOGIC; 
  signal blk00000003_sig0000041b : STD_LOGIC; 
  signal blk00000003_sig0000041a : STD_LOGIC; 
  signal blk00000003_sig00000419 : STD_LOGIC; 
  signal blk00000003_sig00000418 : STD_LOGIC; 
  signal blk00000003_sig00000417 : STD_LOGIC; 
  signal blk00000003_sig00000416 : STD_LOGIC; 
  signal blk00000003_sig00000415 : STD_LOGIC; 
  signal blk00000003_sig00000414 : STD_LOGIC; 
  signal blk00000003_sig00000413 : STD_LOGIC; 
  signal blk00000003_sig00000412 : STD_LOGIC; 
  signal blk00000003_sig00000411 : STD_LOGIC; 
  signal blk00000003_sig00000410 : STD_LOGIC; 
  signal blk00000003_sig0000040f : STD_LOGIC; 
  signal blk00000003_sig0000040e : STD_LOGIC; 
  signal blk00000003_sig0000040d : STD_LOGIC; 
  signal blk00000003_sig0000040c : STD_LOGIC; 
  signal blk00000003_sig0000040b : STD_LOGIC; 
  signal blk00000003_sig0000040a : STD_LOGIC; 
  signal blk00000003_sig00000409 : STD_LOGIC; 
  signal blk00000003_sig00000408 : STD_LOGIC; 
  signal blk00000003_sig00000407 : STD_LOGIC; 
  signal blk00000003_sig00000406 : STD_LOGIC; 
  signal blk00000003_sig00000405 : STD_LOGIC; 
  signal blk00000003_sig00000404 : STD_LOGIC; 
  signal blk00000003_sig00000403 : STD_LOGIC; 
  signal blk00000003_sig00000402 : STD_LOGIC; 
  signal blk00000003_sig00000401 : STD_LOGIC; 
  signal blk00000003_sig00000400 : STD_LOGIC; 
  signal blk00000003_sig000003ff : STD_LOGIC; 
  signal blk00000003_sig000003fe : STD_LOGIC; 
  signal blk00000003_sig000003fd : STD_LOGIC; 
  signal blk00000003_sig000003fc : STD_LOGIC; 
  signal blk00000003_sig000003fb : STD_LOGIC; 
  signal blk00000003_sig000003fa : STD_LOGIC; 
  signal blk00000003_sig000003f9 : STD_LOGIC; 
  signal blk00000003_sig000003f8 : STD_LOGIC; 
  signal blk00000003_sig000003f7 : STD_LOGIC; 
  signal blk00000003_sig000003f6 : STD_LOGIC; 
  signal blk00000003_sig000003f5 : STD_LOGIC; 
  signal blk00000003_sig000003f4 : STD_LOGIC; 
  signal blk00000003_sig000003f3 : STD_LOGIC; 
  signal blk00000003_sig000003f2 : STD_LOGIC; 
  signal blk00000003_sig000003f1 : STD_LOGIC; 
  signal blk00000003_sig000003f0 : STD_LOGIC; 
  signal blk00000003_sig000003ef : STD_LOGIC; 
  signal blk00000003_sig000003ee : STD_LOGIC; 
  signal blk00000003_sig000003ed : STD_LOGIC; 
  signal blk00000003_sig000003ec : STD_LOGIC; 
  signal blk00000003_sig000003eb : STD_LOGIC; 
  signal blk00000003_sig000003ea : STD_LOGIC; 
  signal blk00000003_sig000003e9 : STD_LOGIC; 
  signal blk00000003_sig000003e8 : STD_LOGIC; 
  signal blk00000003_sig000003e7 : STD_LOGIC; 
  signal blk00000003_sig000003e6 : STD_LOGIC; 
  signal blk00000003_sig000003e5 : STD_LOGIC; 
  signal blk00000003_sig000003e4 : STD_LOGIC; 
  signal blk00000003_sig000003e3 : STD_LOGIC; 
  signal blk00000003_sig000003e2 : STD_LOGIC; 
  signal blk00000003_sig000003e1 : STD_LOGIC; 
  signal blk00000003_sig000003e0 : STD_LOGIC; 
  signal blk00000003_sig000003df : STD_LOGIC; 
  signal blk00000003_sig000003de : STD_LOGIC; 
  signal blk00000003_sig000003dd : STD_LOGIC; 
  signal blk00000003_sig000003dc : STD_LOGIC; 
  signal blk00000003_sig000003db : STD_LOGIC; 
  signal blk00000003_sig000003da : STD_LOGIC; 
  signal blk00000003_sig000003d9 : STD_LOGIC; 
  signal blk00000003_sig000003d8 : STD_LOGIC; 
  signal blk00000003_sig000003d7 : STD_LOGIC; 
  signal blk00000003_sig000003d6 : STD_LOGIC; 
  signal blk00000003_sig000003d5 : STD_LOGIC; 
  signal blk00000003_sig000003d4 : STD_LOGIC; 
  signal blk00000003_sig000003d3 : STD_LOGIC; 
  signal blk00000003_sig000003d2 : STD_LOGIC; 
  signal blk00000003_sig000003d1 : STD_LOGIC; 
  signal blk00000003_sig000003d0 : STD_LOGIC; 
  signal blk00000003_sig000003cf : STD_LOGIC; 
  signal blk00000003_sig000003ce : STD_LOGIC; 
  signal blk00000003_sig000003cd : STD_LOGIC; 
  signal blk00000003_sig000003cc : STD_LOGIC; 
  signal blk00000003_sig000003cb : STD_LOGIC; 
  signal blk00000003_sig000003ca : STD_LOGIC; 
  signal blk00000003_sig000003c9 : STD_LOGIC; 
  signal blk00000003_sig000003c8 : STD_LOGIC; 
  signal blk00000003_sig000003c7 : STD_LOGIC; 
  signal blk00000003_sig000003c6 : STD_LOGIC; 
  signal blk00000003_sig000003c5 : STD_LOGIC; 
  signal blk00000003_sig000003c4 : STD_LOGIC; 
  signal blk00000003_sig000003c3 : STD_LOGIC; 
  signal blk00000003_sig000003c2 : STD_LOGIC; 
  signal blk00000003_sig000003c1 : STD_LOGIC; 
  signal blk00000003_sig000003c0 : STD_LOGIC; 
  signal blk00000003_sig000003bf : STD_LOGIC; 
  signal blk00000003_sig000003be : STD_LOGIC; 
  signal blk00000003_sig000003bd : STD_LOGIC; 
  signal blk00000003_sig000003bc : STD_LOGIC; 
  signal blk00000003_sig000003bb : STD_LOGIC; 
  signal blk00000003_sig000003ba : STD_LOGIC; 
  signal blk00000003_sig000003b9 : STD_LOGIC; 
  signal blk00000003_sig000003b8 : STD_LOGIC; 
  signal blk00000003_sig000003b7 : STD_LOGIC; 
  signal blk00000003_sig000003b6 : STD_LOGIC; 
  signal blk00000003_sig000003b5 : STD_LOGIC; 
  signal blk00000003_sig000003b4 : STD_LOGIC; 
  signal blk00000003_sig000003b3 : STD_LOGIC; 
  signal blk00000003_sig000003b2 : STD_LOGIC; 
  signal blk00000003_sig000003b1 : STD_LOGIC; 
  signal blk00000003_sig000003b0 : STD_LOGIC; 
  signal blk00000003_sig000003af : STD_LOGIC; 
  signal blk00000003_sig000003ae : STD_LOGIC; 
  signal blk00000003_sig000003ad : STD_LOGIC; 
  signal blk00000003_sig000003ac : STD_LOGIC; 
  signal blk00000003_sig000003ab : STD_LOGIC; 
  signal blk00000003_sig000003aa : STD_LOGIC; 
  signal blk00000003_sig000003a9 : STD_LOGIC; 
  signal blk00000003_sig000003a8 : STD_LOGIC; 
  signal blk00000003_sig000003a7 : STD_LOGIC; 
  signal blk00000003_sig000003a6 : STD_LOGIC; 
  signal blk00000003_sig000003a5 : STD_LOGIC; 
  signal blk00000003_sig000003a4 : STD_LOGIC; 
  signal blk00000003_sig000003a3 : STD_LOGIC; 
  signal blk00000003_sig000003a2 : STD_LOGIC; 
  signal blk00000003_sig000003a1 : STD_LOGIC; 
  signal blk00000003_sig000003a0 : STD_LOGIC; 
  signal blk00000003_sig0000039f : STD_LOGIC; 
  signal blk00000003_sig0000039e : STD_LOGIC; 
  signal blk00000003_sig0000039d : STD_LOGIC; 
  signal blk00000003_sig0000039c : STD_LOGIC; 
  signal blk00000003_sig0000039b : STD_LOGIC; 
  signal blk00000003_sig0000039a : STD_LOGIC; 
  signal blk00000003_sig00000399 : STD_LOGIC; 
  signal blk00000003_sig00000398 : STD_LOGIC; 
  signal blk00000003_sig00000397 : STD_LOGIC; 
  signal blk00000003_sig00000396 : STD_LOGIC; 
  signal blk00000003_sig00000395 : STD_LOGIC; 
  signal blk00000003_sig00000394 : STD_LOGIC; 
  signal blk00000003_sig00000393 : STD_LOGIC; 
  signal blk00000003_sig00000392 : STD_LOGIC; 
  signal blk00000003_sig00000391 : STD_LOGIC; 
  signal blk00000003_sig00000390 : STD_LOGIC; 
  signal blk00000003_sig0000038f : STD_LOGIC; 
  signal blk00000003_sig0000038e : STD_LOGIC; 
  signal blk00000003_sig0000038d : STD_LOGIC; 
  signal blk00000003_sig0000038c : STD_LOGIC; 
  signal blk00000003_sig0000038b : STD_LOGIC; 
  signal blk00000003_sig0000038a : STD_LOGIC; 
  signal blk00000003_sig00000389 : STD_LOGIC; 
  signal blk00000003_sig00000388 : STD_LOGIC; 
  signal blk00000003_sig00000387 : STD_LOGIC; 
  signal blk00000003_sig00000386 : STD_LOGIC; 
  signal blk00000003_sig00000385 : STD_LOGIC; 
  signal blk00000003_sig00000384 : STD_LOGIC; 
  signal blk00000003_sig00000383 : STD_LOGIC; 
  signal blk00000003_sig00000382 : STD_LOGIC; 
  signal blk00000003_sig00000381 : STD_LOGIC; 
  signal blk00000003_sig00000380 : STD_LOGIC; 
  signal blk00000003_sig0000037f : STD_LOGIC; 
  signal blk00000003_sig0000037e : STD_LOGIC; 
  signal blk00000003_sig0000037d : STD_LOGIC; 
  signal blk00000003_sig0000037c : STD_LOGIC; 
  signal blk00000003_sig0000037b : STD_LOGIC; 
  signal blk00000003_sig0000037a : STD_LOGIC; 
  signal blk00000003_sig00000379 : STD_LOGIC; 
  signal blk00000003_sig00000378 : STD_LOGIC; 
  signal blk00000003_sig00000377 : STD_LOGIC; 
  signal blk00000003_sig00000376 : STD_LOGIC; 
  signal blk00000003_sig00000375 : STD_LOGIC; 
  signal blk00000003_sig00000374 : STD_LOGIC; 
  signal blk00000003_sig00000373 : STD_LOGIC; 
  signal blk00000003_sig00000372 : STD_LOGIC; 
  signal blk00000003_sig00000371 : STD_LOGIC; 
  signal blk00000003_sig00000370 : STD_LOGIC; 
  signal blk00000003_sig0000036f : STD_LOGIC; 
  signal blk00000003_sig0000036e : STD_LOGIC; 
  signal blk00000003_sig0000036d : STD_LOGIC; 
  signal blk00000003_sig0000036c : STD_LOGIC; 
  signal blk00000003_sig0000036b : STD_LOGIC; 
  signal blk00000003_sig0000036a : STD_LOGIC; 
  signal blk00000003_sig00000369 : STD_LOGIC; 
  signal blk00000003_sig00000368 : STD_LOGIC; 
  signal blk00000003_sig00000367 : STD_LOGIC; 
  signal blk00000003_sig00000366 : STD_LOGIC; 
  signal blk00000003_sig00000365 : STD_LOGIC; 
  signal blk00000003_sig00000364 : STD_LOGIC; 
  signal blk00000003_sig00000363 : STD_LOGIC; 
  signal blk00000003_sig00000362 : STD_LOGIC; 
  signal blk00000003_sig00000361 : STD_LOGIC; 
  signal blk00000003_sig00000360 : STD_LOGIC; 
  signal blk00000003_sig0000035f : STD_LOGIC; 
  signal blk00000003_sig0000035e : STD_LOGIC; 
  signal blk00000003_sig0000035d : STD_LOGIC; 
  signal blk00000003_sig0000035c : STD_LOGIC; 
  signal blk00000003_sig0000035b : STD_LOGIC; 
  signal blk00000003_sig0000035a : STD_LOGIC; 
  signal blk00000003_sig00000359 : STD_LOGIC; 
  signal blk00000003_sig00000358 : STD_LOGIC; 
  signal blk00000003_sig00000357 : STD_LOGIC; 
  signal blk00000003_sig00000356 : STD_LOGIC; 
  signal blk00000003_sig00000355 : STD_LOGIC; 
  signal blk00000003_sig00000354 : STD_LOGIC; 
  signal blk00000003_sig00000353 : STD_LOGIC; 
  signal blk00000003_sig00000352 : STD_LOGIC; 
  signal blk00000003_sig00000351 : STD_LOGIC; 
  signal blk00000003_sig00000350 : STD_LOGIC; 
  signal blk00000003_sig0000034f : STD_LOGIC; 
  signal blk00000003_sig0000034e : STD_LOGIC; 
  signal blk00000003_sig0000034d : STD_LOGIC; 
  signal blk00000003_sig0000034c : STD_LOGIC; 
  signal blk00000003_sig0000034b : STD_LOGIC; 
  signal blk00000003_sig0000034a : STD_LOGIC; 
  signal blk00000003_sig00000349 : STD_LOGIC; 
  signal blk00000003_sig00000348 : STD_LOGIC; 
  signal blk00000003_sig00000347 : STD_LOGIC; 
  signal blk00000003_sig00000346 : STD_LOGIC; 
  signal blk00000003_sig00000345 : STD_LOGIC; 
  signal blk00000003_sig00000344 : STD_LOGIC; 
  signal blk00000003_sig00000343 : STD_LOGIC; 
  signal blk00000003_sig00000342 : STD_LOGIC; 
  signal blk00000003_sig00000341 : STD_LOGIC; 
  signal blk00000003_sig00000340 : STD_LOGIC; 
  signal blk00000003_sig0000033f : STD_LOGIC; 
  signal blk00000003_sig0000033e : STD_LOGIC; 
  signal blk00000003_sig0000033d : STD_LOGIC; 
  signal blk00000003_sig0000033c : STD_LOGIC; 
  signal blk00000003_sig0000033b : STD_LOGIC; 
  signal blk00000003_sig0000033a : STD_LOGIC; 
  signal blk00000003_sig00000339 : STD_LOGIC; 
  signal blk00000003_sig00000338 : STD_LOGIC; 
  signal blk00000003_sig00000337 : STD_LOGIC; 
  signal blk00000003_sig00000336 : STD_LOGIC; 
  signal blk00000003_sig00000335 : STD_LOGIC; 
  signal blk00000003_sig00000334 : STD_LOGIC; 
  signal blk00000003_sig00000333 : STD_LOGIC; 
  signal blk00000003_sig00000332 : STD_LOGIC; 
  signal blk00000003_sig00000331 : STD_LOGIC; 
  signal blk00000003_sig00000330 : STD_LOGIC; 
  signal blk00000003_sig0000032f : STD_LOGIC; 
  signal blk00000003_sig0000032e : STD_LOGIC; 
  signal blk00000003_sig0000032d : STD_LOGIC; 
  signal blk00000003_sig0000032c : STD_LOGIC; 
  signal blk00000003_sig0000032b : STD_LOGIC; 
  signal blk00000003_sig0000032a : STD_LOGIC; 
  signal blk00000003_sig00000329 : STD_LOGIC; 
  signal blk00000003_sig00000328 : STD_LOGIC; 
  signal blk00000003_sig00000327 : STD_LOGIC; 
  signal blk00000003_sig00000326 : STD_LOGIC; 
  signal blk00000003_sig00000325 : STD_LOGIC; 
  signal blk00000003_sig00000324 : STD_LOGIC; 
  signal blk00000003_sig00000323 : STD_LOGIC; 
  signal blk00000003_sig00000322 : STD_LOGIC; 
  signal blk00000003_sig00000321 : STD_LOGIC; 
  signal blk00000003_sig00000320 : STD_LOGIC; 
  signal blk00000003_sig0000031f : STD_LOGIC; 
  signal blk00000003_sig0000031e : STD_LOGIC; 
  signal blk00000003_sig0000031d : STD_LOGIC; 
  signal blk00000003_sig0000031c : STD_LOGIC; 
  signal blk00000003_sig0000031b : STD_LOGIC; 
  signal blk00000003_sig0000031a : STD_LOGIC; 
  signal blk00000003_sig00000319 : STD_LOGIC; 
  signal blk00000003_sig00000318 : STD_LOGIC; 
  signal blk00000003_sig00000317 : STD_LOGIC; 
  signal blk00000003_sig00000316 : STD_LOGIC; 
  signal blk00000003_sig00000315 : STD_LOGIC; 
  signal blk00000003_sig00000314 : STD_LOGIC; 
  signal blk00000003_sig00000313 : STD_LOGIC; 
  signal blk00000003_sig00000312 : STD_LOGIC; 
  signal blk00000003_sig00000311 : STD_LOGIC; 
  signal blk00000003_sig00000310 : STD_LOGIC; 
  signal blk00000003_sig0000030f : STD_LOGIC; 
  signal blk00000003_sig0000030e : STD_LOGIC; 
  signal blk00000003_sig0000030d : STD_LOGIC; 
  signal blk00000003_sig0000030c : STD_LOGIC; 
  signal blk00000003_sig0000030b : STD_LOGIC; 
  signal blk00000003_sig0000030a : STD_LOGIC; 
  signal blk00000003_sig00000309 : STD_LOGIC; 
  signal blk00000003_sig00000308 : STD_LOGIC; 
  signal blk00000003_sig00000307 : STD_LOGIC; 
  signal blk00000003_sig00000306 : STD_LOGIC; 
  signal blk00000003_sig00000305 : STD_LOGIC; 
  signal blk00000003_sig00000304 : STD_LOGIC; 
  signal blk00000003_sig00000303 : STD_LOGIC; 
  signal blk00000003_sig00000302 : STD_LOGIC; 
  signal blk00000003_sig00000301 : STD_LOGIC; 
  signal blk00000003_sig00000300 : STD_LOGIC; 
  signal blk00000003_sig000002ff : STD_LOGIC; 
  signal blk00000003_sig000002fe : STD_LOGIC; 
  signal blk00000003_sig000002fd : STD_LOGIC; 
  signal blk00000003_sig000002fc : STD_LOGIC; 
  signal blk00000003_sig000002fb : STD_LOGIC; 
  signal blk00000003_sig000002fa : STD_LOGIC; 
  signal blk00000003_sig000002f9 : STD_LOGIC; 
  signal blk00000003_sig000002f8 : STD_LOGIC; 
  signal blk00000003_sig000002f7 : STD_LOGIC; 
  signal blk00000003_sig000002f6 : STD_LOGIC; 
  signal blk00000003_sig000002f5 : STD_LOGIC; 
  signal blk00000003_sig000002f4 : STD_LOGIC; 
  signal blk00000003_sig000002f3 : STD_LOGIC; 
  signal blk00000003_sig000002f2 : STD_LOGIC; 
  signal blk00000003_sig000002f1 : STD_LOGIC; 
  signal blk00000003_sig000002f0 : STD_LOGIC; 
  signal blk00000003_sig000002ef : STD_LOGIC; 
  signal blk00000003_sig000002ee : STD_LOGIC; 
  signal blk00000003_sig000002ed : STD_LOGIC; 
  signal blk00000003_sig000002ec : STD_LOGIC; 
  signal blk00000003_sig000002eb : STD_LOGIC; 
  signal blk00000003_sig000002ea : STD_LOGIC; 
  signal blk00000003_sig000002e9 : STD_LOGIC; 
  signal blk00000003_sig000002e8 : STD_LOGIC; 
  signal blk00000003_sig000002e7 : STD_LOGIC; 
  signal blk00000003_sig000002e6 : STD_LOGIC; 
  signal blk00000003_sig000002e5 : STD_LOGIC; 
  signal blk00000003_sig000002e4 : STD_LOGIC; 
  signal blk00000003_sig000002e3 : STD_LOGIC; 
  signal blk00000003_sig000002e2 : STD_LOGIC; 
  signal blk00000003_sig000002e1 : STD_LOGIC; 
  signal blk00000003_sig000002e0 : STD_LOGIC; 
  signal blk00000003_sig000002df : STD_LOGIC; 
  signal blk00000003_sig000002de : STD_LOGIC; 
  signal blk00000003_sig000002dd : STD_LOGIC; 
  signal blk00000003_sig000002dc : STD_LOGIC; 
  signal blk00000003_sig000002db : STD_LOGIC; 
  signal blk00000003_sig000002da : STD_LOGIC; 
  signal blk00000003_sig000002d9 : STD_LOGIC; 
  signal blk00000003_sig000002d8 : STD_LOGIC; 
  signal blk00000003_sig000002d7 : STD_LOGIC; 
  signal blk00000003_sig000002d6 : STD_LOGIC; 
  signal blk00000003_sig000002d5 : STD_LOGIC; 
  signal blk00000003_sig000002d4 : STD_LOGIC; 
  signal blk00000003_sig000002d3 : STD_LOGIC; 
  signal blk00000003_sig000002d2 : STD_LOGIC; 
  signal blk00000003_sig000002d1 : STD_LOGIC; 
  signal blk00000003_sig000002d0 : STD_LOGIC; 
  signal blk00000003_sig000002cf : STD_LOGIC; 
  signal blk00000003_sig000002ce : STD_LOGIC; 
  signal blk00000003_sig000002cd : STD_LOGIC; 
  signal blk00000003_sig000002cc : STD_LOGIC; 
  signal blk00000003_sig000002cb : STD_LOGIC; 
  signal blk00000003_sig000002ca : STD_LOGIC; 
  signal blk00000003_sig000002c9 : STD_LOGIC; 
  signal blk00000003_sig000002c8 : STD_LOGIC; 
  signal blk00000003_sig000002c7 : STD_LOGIC; 
  signal blk00000003_sig000002c6 : STD_LOGIC; 
  signal blk00000003_sig000002c5 : STD_LOGIC; 
  signal blk00000003_sig000002c4 : STD_LOGIC; 
  signal blk00000003_sig000002c3 : STD_LOGIC; 
  signal blk00000003_sig000002c2 : STD_LOGIC; 
  signal blk00000003_sig000002c1 : STD_LOGIC; 
  signal blk00000003_sig000002c0 : STD_LOGIC; 
  signal blk00000003_sig000002bf : STD_LOGIC; 
  signal blk00000003_sig000002be : STD_LOGIC; 
  signal blk00000003_sig000002bd : STD_LOGIC; 
  signal blk00000003_sig000002bc : STD_LOGIC; 
  signal blk00000003_sig000002bb : STD_LOGIC; 
  signal blk00000003_sig000002ba : STD_LOGIC; 
  signal blk00000003_sig000002b9 : STD_LOGIC; 
  signal blk00000003_sig000002b8 : STD_LOGIC; 
  signal blk00000003_sig000002b7 : STD_LOGIC; 
  signal blk00000003_sig000002b6 : STD_LOGIC; 
  signal blk00000003_sig000002b5 : STD_LOGIC; 
  signal blk00000003_sig000002b4 : STD_LOGIC; 
  signal blk00000003_sig000002b3 : STD_LOGIC; 
  signal blk00000003_sig000002b2 : STD_LOGIC; 
  signal blk00000003_sig000002b1 : STD_LOGIC; 
  signal blk00000003_sig000002b0 : STD_LOGIC; 
  signal blk00000003_sig000002af : STD_LOGIC; 
  signal blk00000003_sig000002ae : STD_LOGIC; 
  signal blk00000003_sig000002ad : STD_LOGIC; 
  signal blk00000003_sig000002ac : STD_LOGIC; 
  signal blk00000003_sig000002ab : STD_LOGIC; 
  signal blk00000003_sig000002aa : STD_LOGIC; 
  signal blk00000003_sig000002a9 : STD_LOGIC; 
  signal blk00000003_sig000002a8 : STD_LOGIC; 
  signal blk00000003_sig000002a7 : STD_LOGIC; 
  signal blk00000003_sig000002a6 : STD_LOGIC; 
  signal blk00000003_sig000002a5 : STD_LOGIC; 
  signal blk00000003_sig000002a4 : STD_LOGIC; 
  signal blk00000003_sig000002a3 : STD_LOGIC; 
  signal blk00000003_sig000002a2 : STD_LOGIC; 
  signal blk00000003_sig000002a1 : STD_LOGIC; 
  signal blk00000003_sig000002a0 : STD_LOGIC; 
  signal blk00000003_sig0000029f : STD_LOGIC; 
  signal blk00000003_sig0000029e : STD_LOGIC; 
  signal blk00000003_sig0000029d : STD_LOGIC; 
  signal blk00000003_sig0000029c : STD_LOGIC; 
  signal blk00000003_sig0000029b : STD_LOGIC; 
  signal blk00000003_sig0000029a : STD_LOGIC; 
  signal blk00000003_sig00000299 : STD_LOGIC; 
  signal blk00000003_sig00000298 : STD_LOGIC; 
  signal blk00000003_sig00000297 : STD_LOGIC; 
  signal blk00000003_sig00000296 : STD_LOGIC; 
  signal blk00000003_sig00000295 : STD_LOGIC; 
  signal blk00000003_sig00000294 : STD_LOGIC; 
  signal blk00000003_sig00000293 : STD_LOGIC; 
  signal blk00000003_sig00000292 : STD_LOGIC; 
  signal blk00000003_sig00000291 : STD_LOGIC; 
  signal blk00000003_sig00000290 : STD_LOGIC; 
  signal blk00000003_sig0000028f : STD_LOGIC; 
  signal blk00000003_sig0000028e : STD_LOGIC; 
  signal blk00000003_sig0000028d : STD_LOGIC; 
  signal blk00000003_sig0000028c : STD_LOGIC; 
  signal blk00000003_sig0000028b : STD_LOGIC; 
  signal blk00000003_sig0000028a : STD_LOGIC; 
  signal blk00000003_sig00000289 : STD_LOGIC; 
  signal blk00000003_sig00000288 : STD_LOGIC; 
  signal blk00000003_sig00000287 : STD_LOGIC; 
  signal blk00000003_sig00000286 : STD_LOGIC; 
  signal blk00000003_sig00000285 : STD_LOGIC; 
  signal blk00000003_sig00000284 : STD_LOGIC; 
  signal blk00000003_sig00000283 : STD_LOGIC; 
  signal blk00000003_sig00000282 : STD_LOGIC; 
  signal blk00000003_sig00000281 : STD_LOGIC; 
  signal blk00000003_sig00000280 : STD_LOGIC; 
  signal blk00000003_sig0000027f : STD_LOGIC; 
  signal blk00000003_sig0000027e : STD_LOGIC; 
  signal blk00000003_sig0000027d : STD_LOGIC; 
  signal blk00000003_sig0000027c : STD_LOGIC; 
  signal blk00000003_sig0000027b : STD_LOGIC; 
  signal blk00000003_sig0000027a : STD_LOGIC; 
  signal blk00000003_sig00000279 : STD_LOGIC; 
  signal blk00000003_sig00000278 : STD_LOGIC; 
  signal blk00000003_sig00000277 : STD_LOGIC; 
  signal blk00000003_sig00000276 : STD_LOGIC; 
  signal blk00000003_sig00000275 : STD_LOGIC; 
  signal blk00000003_sig00000274 : STD_LOGIC; 
  signal blk00000003_sig00000273 : STD_LOGIC; 
  signal blk00000003_sig00000272 : STD_LOGIC; 
  signal blk00000003_sig00000271 : STD_LOGIC; 
  signal blk00000003_sig00000270 : STD_LOGIC; 
  signal blk00000003_sig0000026f : STD_LOGIC; 
  signal blk00000003_sig0000026e : STD_LOGIC; 
  signal blk00000003_sig0000026d : STD_LOGIC; 
  signal blk00000003_sig0000026c : STD_LOGIC; 
  signal blk00000003_sig0000026b : STD_LOGIC; 
  signal blk00000003_sig0000026a : STD_LOGIC; 
  signal blk00000003_sig00000269 : STD_LOGIC; 
  signal blk00000003_sig00000268 : STD_LOGIC; 
  signal blk00000003_sig00000267 : STD_LOGIC; 
  signal blk00000003_sig00000266 : STD_LOGIC; 
  signal blk00000003_sig00000265 : STD_LOGIC; 
  signal blk00000003_sig00000264 : STD_LOGIC; 
  signal blk00000003_sig00000263 : STD_LOGIC; 
  signal blk00000003_sig00000262 : STD_LOGIC; 
  signal blk00000003_sig00000261 : STD_LOGIC; 
  signal blk00000003_sig00000260 : STD_LOGIC; 
  signal blk00000003_sig0000025f : STD_LOGIC; 
  signal blk00000003_sig0000025e : STD_LOGIC; 
  signal blk00000003_sig0000025d : STD_LOGIC; 
  signal blk00000003_sig0000025c : STD_LOGIC; 
  signal blk00000003_sig0000025b : STD_LOGIC; 
  signal blk00000003_sig0000025a : STD_LOGIC; 
  signal blk00000003_sig00000259 : STD_LOGIC; 
  signal blk00000003_sig00000258 : STD_LOGIC; 
  signal blk00000003_sig00000257 : STD_LOGIC; 
  signal blk00000003_sig00000256 : STD_LOGIC; 
  signal blk00000003_sig00000255 : STD_LOGIC; 
  signal blk00000003_sig00000254 : STD_LOGIC; 
  signal blk00000003_sig00000253 : STD_LOGIC; 
  signal blk00000003_sig00000252 : STD_LOGIC; 
  signal blk00000003_sig00000251 : STD_LOGIC; 
  signal blk00000003_sig00000250 : STD_LOGIC; 
  signal blk00000003_sig0000024f : STD_LOGIC; 
  signal blk00000003_sig0000024e : STD_LOGIC; 
  signal blk00000003_sig0000024d : STD_LOGIC; 
  signal blk00000003_sig0000024c : STD_LOGIC; 
  signal blk00000003_sig0000024b : STD_LOGIC; 
  signal blk00000003_sig0000024a : STD_LOGIC; 
  signal blk00000003_sig00000249 : STD_LOGIC; 
  signal blk00000003_sig00000248 : STD_LOGIC; 
  signal blk00000003_sig00000247 : STD_LOGIC; 
  signal blk00000003_sig00000246 : STD_LOGIC; 
  signal blk00000003_sig00000245 : STD_LOGIC; 
  signal blk00000003_sig00000244 : STD_LOGIC; 
  signal blk00000003_sig00000243 : STD_LOGIC; 
  signal blk00000003_sig00000242 : STD_LOGIC; 
  signal blk00000003_sig00000241 : STD_LOGIC; 
  signal blk00000003_sig00000240 : STD_LOGIC; 
  signal blk00000003_sig0000023f : STD_LOGIC; 
  signal blk00000003_sig0000023e : STD_LOGIC; 
  signal blk00000003_sig0000023d : STD_LOGIC; 
  signal blk00000003_sig0000023c : STD_LOGIC; 
  signal blk00000003_sig0000023b : STD_LOGIC; 
  signal blk00000003_sig0000023a : STD_LOGIC; 
  signal blk00000003_sig00000239 : STD_LOGIC; 
  signal blk00000003_sig00000238 : STD_LOGIC; 
  signal blk00000003_sig00000237 : STD_LOGIC; 
  signal blk00000003_sig00000236 : STD_LOGIC; 
  signal blk00000003_sig00000235 : STD_LOGIC; 
  signal blk00000003_sig00000234 : STD_LOGIC; 
  signal blk00000003_sig00000233 : STD_LOGIC; 
  signal blk00000003_sig00000232 : STD_LOGIC; 
  signal blk00000003_sig00000231 : STD_LOGIC; 
  signal blk00000003_sig00000230 : STD_LOGIC; 
  signal blk00000003_sig0000022f : STD_LOGIC; 
  signal blk00000003_sig0000022e : STD_LOGIC; 
  signal blk00000003_sig0000022d : STD_LOGIC; 
  signal blk00000003_sig0000022c : STD_LOGIC; 
  signal blk00000003_sig0000022b : STD_LOGIC; 
  signal blk00000003_sig0000022a : STD_LOGIC; 
  signal blk00000003_sig00000229 : STD_LOGIC; 
  signal blk00000003_sig00000228 : STD_LOGIC; 
  signal blk00000003_sig00000227 : STD_LOGIC; 
  signal blk00000003_sig00000226 : STD_LOGIC; 
  signal blk00000003_sig00000225 : STD_LOGIC; 
  signal blk00000003_sig00000224 : STD_LOGIC; 
  signal blk00000003_sig00000223 : STD_LOGIC; 
  signal blk00000003_sig00000222 : STD_LOGIC; 
  signal blk00000003_sig00000221 : STD_LOGIC; 
  signal blk00000003_sig00000220 : STD_LOGIC; 
  signal blk00000003_sig0000021f : STD_LOGIC; 
  signal blk00000003_sig0000021e : STD_LOGIC; 
  signal blk00000003_sig0000021d : STD_LOGIC; 
  signal blk00000003_sig0000021c : STD_LOGIC; 
  signal blk00000003_sig0000021b : STD_LOGIC; 
  signal blk00000003_sig0000021a : STD_LOGIC; 
  signal blk00000003_sig00000219 : STD_LOGIC; 
  signal blk00000003_sig00000218 : STD_LOGIC; 
  signal blk00000003_sig00000217 : STD_LOGIC; 
  signal blk00000003_sig00000216 : STD_LOGIC; 
  signal blk00000003_sig00000215 : STD_LOGIC; 
  signal blk00000003_sig00000214 : STD_LOGIC; 
  signal blk00000003_sig00000213 : STD_LOGIC; 
  signal blk00000003_sig00000212 : STD_LOGIC; 
  signal blk00000003_sig00000211 : STD_LOGIC; 
  signal blk00000003_sig00000210 : STD_LOGIC; 
  signal blk00000003_sig0000020f : STD_LOGIC; 
  signal blk00000003_sig0000020e : STD_LOGIC; 
  signal blk00000003_sig0000020d : STD_LOGIC; 
  signal blk00000003_sig0000020c : STD_LOGIC; 
  signal blk00000003_sig0000020b : STD_LOGIC; 
  signal blk00000003_sig0000020a : STD_LOGIC; 
  signal blk00000003_sig00000209 : STD_LOGIC; 
  signal blk00000003_sig00000208 : STD_LOGIC; 
  signal blk00000003_sig00000207 : STD_LOGIC; 
  signal blk00000003_sig00000206 : STD_LOGIC; 
  signal blk00000003_sig00000205 : STD_LOGIC; 
  signal blk00000003_sig00000204 : STD_LOGIC; 
  signal blk00000003_sig00000203 : STD_LOGIC; 
  signal blk00000003_sig00000202 : STD_LOGIC; 
  signal blk00000003_sig00000201 : STD_LOGIC; 
  signal blk00000003_sig00000200 : STD_LOGIC; 
  signal blk00000003_sig000001ff : STD_LOGIC; 
  signal blk00000003_sig000001fe : STD_LOGIC; 
  signal blk00000003_sig000001fd : STD_LOGIC; 
  signal blk00000003_sig000001fc : STD_LOGIC; 
  signal blk00000003_sig000001fb : STD_LOGIC; 
  signal blk00000003_sig000001fa : STD_LOGIC; 
  signal blk00000003_sig000001f9 : STD_LOGIC; 
  signal blk00000003_sig000001f8 : STD_LOGIC; 
  signal blk00000003_sig000001f7 : STD_LOGIC; 
  signal blk00000003_sig000001f6 : STD_LOGIC; 
  signal blk00000003_sig000001f5 : STD_LOGIC; 
  signal blk00000003_sig000001f4 : STD_LOGIC; 
  signal blk00000003_sig000001f3 : STD_LOGIC; 
  signal blk00000003_sig000001f2 : STD_LOGIC; 
  signal blk00000003_sig000001f1 : STD_LOGIC; 
  signal blk00000003_sig000001f0 : STD_LOGIC; 
  signal blk00000003_sig000001ef : STD_LOGIC; 
  signal blk00000003_sig000001ee : STD_LOGIC; 
  signal blk00000003_sig000001ed : STD_LOGIC; 
  signal blk00000003_sig000001ec : STD_LOGIC; 
  signal blk00000003_sig000001eb : STD_LOGIC; 
  signal blk00000003_sig000001ea : STD_LOGIC; 
  signal blk00000003_sig000001e9 : STD_LOGIC; 
  signal blk00000003_sig000001e8 : STD_LOGIC; 
  signal blk00000003_sig000001e7 : STD_LOGIC; 
  signal blk00000003_sig000001e6 : STD_LOGIC; 
  signal blk00000003_sig000001e5 : STD_LOGIC; 
  signal blk00000003_sig000001e4 : STD_LOGIC; 
  signal blk00000003_sig000001e3 : STD_LOGIC; 
  signal blk00000003_sig000001e2 : STD_LOGIC; 
  signal blk00000003_sig000001e1 : STD_LOGIC; 
  signal blk00000003_sig000001e0 : STD_LOGIC; 
  signal blk00000003_sig000001df : STD_LOGIC; 
  signal blk00000003_sig000001de : STD_LOGIC; 
  signal blk00000003_sig000001dd : STD_LOGIC; 
  signal blk00000003_sig000001dc : STD_LOGIC; 
  signal blk00000003_sig000001db : STD_LOGIC; 
  signal blk00000003_sig000001da : STD_LOGIC; 
  signal blk00000003_sig000001d9 : STD_LOGIC; 
  signal blk00000003_sig000001d8 : STD_LOGIC; 
  signal blk00000003_sig000001d7 : STD_LOGIC; 
  signal blk00000003_sig000001d6 : STD_LOGIC; 
  signal blk00000003_sig000001d5 : STD_LOGIC; 
  signal blk00000003_sig000001d4 : STD_LOGIC; 
  signal blk00000003_sig000001d3 : STD_LOGIC; 
  signal blk00000003_sig000001d2 : STD_LOGIC; 
  signal blk00000003_sig000001d1 : STD_LOGIC; 
  signal blk00000003_sig000001d0 : STD_LOGIC; 
  signal blk00000003_sig000001cf : STD_LOGIC; 
  signal blk00000003_sig000001ce : STD_LOGIC; 
  signal blk00000003_sig000001cd : STD_LOGIC; 
  signal blk00000003_sig000001cc : STD_LOGIC; 
  signal blk00000003_sig000001cb : STD_LOGIC; 
  signal blk00000003_sig000001ca : STD_LOGIC; 
  signal blk00000003_sig000001c9 : STD_LOGIC; 
  signal blk00000003_sig000001c8 : STD_LOGIC; 
  signal blk00000003_sig000001c7 : STD_LOGIC; 
  signal blk00000003_sig000001c6 : STD_LOGIC; 
  signal blk00000003_sig000001c5 : STD_LOGIC; 
  signal blk00000003_sig000001c4 : STD_LOGIC; 
  signal blk00000003_sig000001c3 : STD_LOGIC; 
  signal blk00000003_sig000001c2 : STD_LOGIC; 
  signal blk00000003_sig000001c1 : STD_LOGIC; 
  signal blk00000003_sig000001c0 : STD_LOGIC; 
  signal blk00000003_sig000001bf : STD_LOGIC; 
  signal blk00000003_sig000001be : STD_LOGIC; 
  signal blk00000003_sig000001bd : STD_LOGIC; 
  signal blk00000003_sig000001bc : STD_LOGIC; 
  signal blk00000003_sig000001bb : STD_LOGIC; 
  signal blk00000003_sig000001ba : STD_LOGIC; 
  signal blk00000003_sig000001b9 : STD_LOGIC; 
  signal blk00000003_sig000001b8 : STD_LOGIC; 
  signal blk00000003_sig000001b7 : STD_LOGIC; 
  signal blk00000003_sig000001b6 : STD_LOGIC; 
  signal blk00000003_sig000001b5 : STD_LOGIC; 
  signal blk00000003_sig000001b4 : STD_LOGIC; 
  signal blk00000003_sig000001b3 : STD_LOGIC; 
  signal blk00000003_sig000001b2 : STD_LOGIC; 
  signal blk00000003_sig000001b1 : STD_LOGIC; 
  signal blk00000003_sig000001b0 : STD_LOGIC; 
  signal blk00000003_sig000001af : STD_LOGIC; 
  signal blk00000003_sig000001ae : STD_LOGIC; 
  signal blk00000003_sig000001ad : STD_LOGIC; 
  signal blk00000003_sig000001ac : STD_LOGIC; 
  signal blk00000003_sig000001ab : STD_LOGIC; 
  signal blk00000003_sig000001aa : STD_LOGIC; 
  signal blk00000003_sig000001a9 : STD_LOGIC; 
  signal blk00000003_sig000001a8 : STD_LOGIC; 
  signal blk00000003_sig000001a7 : STD_LOGIC; 
  signal blk00000003_sig000001a6 : STD_LOGIC; 
  signal blk00000003_sig000001a5 : STD_LOGIC; 
  signal blk00000003_sig000001a4 : STD_LOGIC; 
  signal blk00000003_sig000001a3 : STD_LOGIC; 
  signal blk00000003_sig000001a2 : STD_LOGIC; 
  signal blk00000003_sig000001a1 : STD_LOGIC; 
  signal blk00000003_sig000001a0 : STD_LOGIC; 
  signal blk00000003_sig0000019f : STD_LOGIC; 
  signal blk00000003_sig0000019e : STD_LOGIC; 
  signal blk00000003_sig0000019d : STD_LOGIC; 
  signal blk00000003_sig0000019c : STD_LOGIC; 
  signal blk00000003_sig0000019b : STD_LOGIC; 
  signal blk00000003_sig0000019a : STD_LOGIC; 
  signal blk00000003_sig00000199 : STD_LOGIC; 
  signal blk00000003_sig00000198 : STD_LOGIC; 
  signal blk00000003_sig00000197 : STD_LOGIC; 
  signal blk00000003_sig00000196 : STD_LOGIC; 
  signal blk00000003_sig00000195 : STD_LOGIC; 
  signal blk00000003_sig00000194 : STD_LOGIC; 
  signal blk00000003_sig00000193 : STD_LOGIC; 
  signal blk00000003_sig00000192 : STD_LOGIC; 
  signal blk00000003_sig00000191 : STD_LOGIC; 
  signal blk00000003_sig00000190 : STD_LOGIC; 
  signal blk00000003_sig0000018f : STD_LOGIC; 
  signal blk00000003_sig0000018e : STD_LOGIC; 
  signal blk00000003_sig0000018d : STD_LOGIC; 
  signal blk00000003_sig0000018c : STD_LOGIC; 
  signal blk00000003_sig0000018b : STD_LOGIC; 
  signal blk00000003_sig0000018a : STD_LOGIC; 
  signal blk00000003_sig00000189 : STD_LOGIC; 
  signal blk00000003_sig00000188 : STD_LOGIC; 
  signal blk00000003_sig00000187 : STD_LOGIC; 
  signal blk00000003_sig00000186 : STD_LOGIC; 
  signal blk00000003_sig00000185 : STD_LOGIC; 
  signal blk00000003_sig00000184 : STD_LOGIC; 
  signal blk00000003_sig00000183 : STD_LOGIC; 
  signal blk00000003_sig00000182 : STD_LOGIC; 
  signal blk00000003_sig00000181 : STD_LOGIC; 
  signal blk00000003_sig00000180 : STD_LOGIC; 
  signal blk00000003_sig0000017f : STD_LOGIC; 
  signal blk00000003_sig0000017e : STD_LOGIC; 
  signal blk00000003_sig0000017d : STD_LOGIC; 
  signal blk00000003_sig0000017c : STD_LOGIC; 
  signal blk00000003_sig0000017b : STD_LOGIC; 
  signal blk00000003_sig0000017a : STD_LOGIC; 
  signal blk00000003_sig00000179 : STD_LOGIC; 
  signal blk00000003_sig00000178 : STD_LOGIC; 
  signal blk00000003_sig00000177 : STD_LOGIC; 
  signal blk00000003_sig00000176 : STD_LOGIC; 
  signal blk00000003_sig00000175 : STD_LOGIC; 
  signal blk00000003_sig00000174 : STD_LOGIC; 
  signal blk00000003_sig00000173 : STD_LOGIC; 
  signal blk00000003_sig00000172 : STD_LOGIC; 
  signal blk00000003_sig00000171 : STD_LOGIC; 
  signal blk00000003_sig00000170 : STD_LOGIC; 
  signal blk00000003_sig0000016f : STD_LOGIC; 
  signal blk00000003_sig0000016e : STD_LOGIC; 
  signal blk00000003_sig0000016d : STD_LOGIC; 
  signal blk00000003_sig0000016c : STD_LOGIC; 
  signal blk00000003_sig0000016b : STD_LOGIC; 
  signal blk00000003_sig0000016a : STD_LOGIC; 
  signal blk00000003_sig00000169 : STD_LOGIC; 
  signal blk00000003_sig00000168 : STD_LOGIC; 
  signal blk00000003_sig00000167 : STD_LOGIC; 
  signal blk00000003_sig00000166 : STD_LOGIC; 
  signal blk00000003_sig00000165 : STD_LOGIC; 
  signal blk00000003_sig00000164 : STD_LOGIC; 
  signal blk00000003_sig00000163 : STD_LOGIC; 
  signal blk00000003_sig00000162 : STD_LOGIC; 
  signal blk00000003_sig00000161 : STD_LOGIC; 
  signal blk00000003_sig00000160 : STD_LOGIC; 
  signal blk00000003_sig0000015f : STD_LOGIC; 
  signal blk00000003_sig0000015e : STD_LOGIC; 
  signal blk00000003_sig0000015d : STD_LOGIC; 
  signal blk00000003_sig0000015c : STD_LOGIC; 
  signal blk00000003_sig0000015b : STD_LOGIC; 
  signal blk00000003_sig0000015a : STD_LOGIC; 
  signal blk00000003_sig00000159 : STD_LOGIC; 
  signal blk00000003_sig00000158 : STD_LOGIC; 
  signal blk00000003_sig00000157 : STD_LOGIC; 
  signal blk00000003_sig00000156 : STD_LOGIC; 
  signal blk00000003_sig00000155 : STD_LOGIC; 
  signal blk00000003_sig00000154 : STD_LOGIC; 
  signal blk00000003_sig00000153 : STD_LOGIC; 
  signal blk00000003_sig00000152 : STD_LOGIC; 
  signal blk00000003_sig00000151 : STD_LOGIC; 
  signal blk00000003_sig00000150 : STD_LOGIC; 
  signal blk00000003_sig0000014f : STD_LOGIC; 
  signal blk00000003_sig0000014e : STD_LOGIC; 
  signal blk00000003_sig0000014d : STD_LOGIC; 
  signal blk00000003_sig0000014c : STD_LOGIC; 
  signal blk00000003_sig0000014b : STD_LOGIC; 
  signal blk00000003_sig0000014a : STD_LOGIC; 
  signal blk00000003_sig00000149 : STD_LOGIC; 
  signal blk00000003_sig00000148 : STD_LOGIC; 
  signal blk00000003_sig00000147 : STD_LOGIC; 
  signal blk00000003_sig00000146 : STD_LOGIC; 
  signal blk00000003_sig00000145 : STD_LOGIC; 
  signal blk00000003_sig00000144 : STD_LOGIC; 
  signal blk00000003_sig00000143 : STD_LOGIC; 
  signal blk00000003_sig00000142 : STD_LOGIC; 
  signal blk00000003_sig00000141 : STD_LOGIC; 
  signal blk00000003_sig00000140 : STD_LOGIC; 
  signal blk00000003_sig0000013f : STD_LOGIC; 
  signal blk00000003_sig0000013e : STD_LOGIC; 
  signal blk00000003_sig0000013d : STD_LOGIC; 
  signal blk00000003_sig0000013c : STD_LOGIC; 
  signal blk00000003_sig0000013b : STD_LOGIC; 
  signal blk00000003_sig0000013a : STD_LOGIC; 
  signal blk00000003_sig00000139 : STD_LOGIC; 
  signal blk00000003_sig00000138 : STD_LOGIC; 
  signal blk00000003_sig00000137 : STD_LOGIC; 
  signal blk00000003_sig00000136 : STD_LOGIC; 
  signal blk00000003_sig00000135 : STD_LOGIC; 
  signal blk00000003_sig00000134 : STD_LOGIC; 
  signal blk00000003_sig00000133 : STD_LOGIC; 
  signal blk00000003_sig00000132 : STD_LOGIC; 
  signal blk00000003_sig00000131 : STD_LOGIC; 
  signal blk00000003_sig00000130 : STD_LOGIC; 
  signal blk00000003_sig0000012f : STD_LOGIC; 
  signal blk00000003_sig0000012e : STD_LOGIC; 
  signal blk00000003_sig0000012d : STD_LOGIC; 
  signal blk00000003_sig0000012c : STD_LOGIC; 
  signal blk00000003_sig0000012b : STD_LOGIC; 
  signal blk00000003_sig0000012a : STD_LOGIC; 
  signal blk00000003_sig00000129 : STD_LOGIC; 
  signal blk00000003_sig00000128 : STD_LOGIC; 
  signal blk00000003_sig00000127 : STD_LOGIC; 
  signal blk00000003_sig00000126 : STD_LOGIC; 
  signal blk00000003_sig00000125 : STD_LOGIC; 
  signal blk00000003_sig00000124 : STD_LOGIC; 
  signal blk00000003_sig00000123 : STD_LOGIC; 
  signal blk00000003_sig00000122 : STD_LOGIC; 
  signal blk00000003_sig00000121 : STD_LOGIC; 
  signal blk00000003_sig00000120 : STD_LOGIC; 
  signal blk00000003_sig0000011f : STD_LOGIC; 
  signal blk00000003_sig0000011e : STD_LOGIC; 
  signal blk00000003_sig0000011d : STD_LOGIC; 
  signal blk00000003_sig0000011c : STD_LOGIC; 
  signal blk00000003_sig0000011b : STD_LOGIC; 
  signal blk00000003_sig0000011a : STD_LOGIC; 
  signal blk00000003_sig00000119 : STD_LOGIC; 
  signal blk00000003_sig00000118 : STD_LOGIC; 
  signal blk00000003_sig00000117 : STD_LOGIC; 
  signal blk00000003_sig00000116 : STD_LOGIC; 
  signal blk00000003_sig00000115 : STD_LOGIC; 
  signal blk00000003_sig00000114 : STD_LOGIC; 
  signal blk00000003_sig00000113 : STD_LOGIC; 
  signal blk00000003_sig00000112 : STD_LOGIC; 
  signal blk00000003_sig00000111 : STD_LOGIC; 
  signal blk00000003_sig00000110 : STD_LOGIC; 
  signal blk00000003_sig0000010f : STD_LOGIC; 
  signal blk00000003_sig0000010e : STD_LOGIC; 
  signal blk00000003_sig0000010d : STD_LOGIC; 
  signal blk00000003_sig0000010c : STD_LOGIC; 
  signal blk00000003_sig0000010b : STD_LOGIC; 
  signal blk00000003_sig0000010a : STD_LOGIC; 
  signal blk00000003_sig00000109 : STD_LOGIC; 
  signal blk00000003_sig00000108 : STD_LOGIC; 
  signal blk00000003_sig00000107 : STD_LOGIC; 
  signal blk00000003_sig00000106 : STD_LOGIC; 
  signal blk00000003_sig00000105 : STD_LOGIC; 
  signal blk00000003_sig00000104 : STD_LOGIC; 
  signal blk00000003_sig00000103 : STD_LOGIC; 
  signal blk00000003_sig00000102 : STD_LOGIC; 
  signal blk00000003_sig00000101 : STD_LOGIC; 
  signal blk00000003_sig00000100 : STD_LOGIC; 
  signal blk00000003_sig000000ff : STD_LOGIC; 
  signal blk00000003_sig000000fe : STD_LOGIC; 
  signal blk00000003_sig000000fd : STD_LOGIC; 
  signal blk00000003_sig000000fc : STD_LOGIC; 
  signal blk00000003_sig000000fb : STD_LOGIC; 
  signal blk00000003_sig000000fa : STD_LOGIC; 
  signal blk00000003_sig000000f9 : STD_LOGIC; 
  signal blk00000003_sig000000f8 : STD_LOGIC; 
  signal blk00000003_sig000000f7 : STD_LOGIC; 
  signal blk00000003_sig000000f6 : STD_LOGIC; 
  signal blk00000003_sig000000f5 : STD_LOGIC; 
  signal blk00000003_sig000000f4 : STD_LOGIC; 
  signal blk00000003_sig000000f3 : STD_LOGIC; 
  signal blk00000003_sig000000f2 : STD_LOGIC; 
  signal blk00000003_sig000000f1 : STD_LOGIC; 
  signal blk00000003_sig000000f0 : STD_LOGIC; 
  signal blk00000003_sig000000ef : STD_LOGIC; 
  signal blk00000003_sig000000ee : STD_LOGIC; 
  signal blk00000003_sig000000ed : STD_LOGIC; 
  signal blk00000003_sig000000ec : STD_LOGIC; 
  signal blk00000003_sig000000eb : STD_LOGIC; 
  signal blk00000003_sig000000ea : STD_LOGIC; 
  signal blk00000003_sig000000e9 : STD_LOGIC; 
  signal blk00000003_sig000000e8 : STD_LOGIC; 
  signal blk00000003_sig000000e7 : STD_LOGIC; 
  signal blk00000003_sig000000e6 : STD_LOGIC; 
  signal blk00000003_sig000000e5 : STD_LOGIC; 
  signal blk00000003_sig000000e4 : STD_LOGIC; 
  signal blk00000003_sig000000e3 : STD_LOGIC; 
  signal blk00000003_sig000000e2 : STD_LOGIC; 
  signal blk00000003_sig000000e1 : STD_LOGIC; 
  signal blk00000003_sig000000e0 : STD_LOGIC; 
  signal blk00000003_sig000000df : STD_LOGIC; 
  signal blk00000003_sig000000de : STD_LOGIC; 
  signal blk00000003_sig000000dd : STD_LOGIC; 
  signal blk00000003_sig000000dc : STD_LOGIC; 
  signal blk00000003_sig000000db : STD_LOGIC; 
  signal blk00000003_sig000000da : STD_LOGIC; 
  signal blk00000003_sig000000d9 : STD_LOGIC; 
  signal blk00000003_sig000000d8 : STD_LOGIC; 
  signal blk00000003_sig000000d7 : STD_LOGIC; 
  signal blk00000003_sig000000d6 : STD_LOGIC; 
  signal blk00000003_sig000000d5 : STD_LOGIC; 
  signal blk00000003_sig000000d4 : STD_LOGIC; 
  signal blk00000003_sig000000d3 : STD_LOGIC; 
  signal blk00000003_sig000000d2 : STD_LOGIC; 
  signal blk00000003_sig000000d1 : STD_LOGIC; 
  signal blk00000003_sig000000d0 : STD_LOGIC; 
  signal blk00000003_sig000000cf : STD_LOGIC; 
  signal blk00000003_sig000000ce : STD_LOGIC; 
  signal blk00000003_sig000000cd : STD_LOGIC; 
  signal blk00000003_sig000000cc : STD_LOGIC; 
  signal blk00000003_sig000000cb : STD_LOGIC; 
  signal blk00000003_sig000000ca : STD_LOGIC; 
  signal blk00000003_sig000000c9 : STD_LOGIC; 
  signal blk00000003_sig000000c8 : STD_LOGIC; 
  signal blk00000003_sig000000c7 : STD_LOGIC; 
  signal blk00000003_sig000000c6 : STD_LOGIC; 
  signal blk00000003_sig000000c5 : STD_LOGIC; 
  signal blk00000003_sig000000c4 : STD_LOGIC; 
  signal blk00000003_sig000000c3 : STD_LOGIC; 
  signal blk00000003_sig000000c2 : STD_LOGIC; 
  signal blk00000003_sig000000c1 : STD_LOGIC; 
  signal blk00000003_sig000000c0 : STD_LOGIC; 
  signal blk00000003_sig000000bf : STD_LOGIC; 
  signal blk00000003_sig000000be : STD_LOGIC; 
  signal blk00000003_sig000000bd : STD_LOGIC; 
  signal blk00000003_sig000000bc : STD_LOGIC; 
  signal blk00000003_sig000000bb : STD_LOGIC; 
  signal blk00000003_sig000000ba : STD_LOGIC; 
  signal blk00000003_sig000000b9 : STD_LOGIC; 
  signal blk00000003_sig000000b8 : STD_LOGIC; 
  signal blk00000003_sig000000b7 : STD_LOGIC; 
  signal blk00000003_sig000000b6 : STD_LOGIC; 
  signal blk00000003_sig000000b5 : STD_LOGIC; 
  signal blk00000003_sig000000b4 : STD_LOGIC; 
  signal blk00000003_sig000000b3 : STD_LOGIC; 
  signal blk00000003_sig000000b2 : STD_LOGIC; 
  signal blk00000003_sig000000b1 : STD_LOGIC; 
  signal blk00000003_sig000000b0 : STD_LOGIC; 
  signal blk00000003_sig000000af : STD_LOGIC; 
  signal blk00000003_sig000000ae : STD_LOGIC; 
  signal blk00000003_sig000000ad : STD_LOGIC; 
  signal blk00000003_sig000000ac : STD_LOGIC; 
  signal blk00000003_sig000000ab : STD_LOGIC; 
  signal blk00000003_sig000000aa : STD_LOGIC; 
  signal blk00000003_sig000000a9 : STD_LOGIC; 
  signal blk00000003_sig000000a8 : STD_LOGIC; 
  signal blk00000003_sig000000a7 : STD_LOGIC; 
  signal blk00000003_sig000000a6 : STD_LOGIC; 
  signal blk00000003_sig000000a5 : STD_LOGIC; 
  signal blk00000003_sig000000a4 : STD_LOGIC; 
  signal blk00000003_sig000000a3 : STD_LOGIC; 
  signal blk00000003_sig000000a2 : STD_LOGIC; 
  signal blk00000003_sig000000a1 : STD_LOGIC; 
  signal blk00000003_sig000000a0 : STD_LOGIC; 
  signal blk00000003_sig0000009f : STD_LOGIC; 
  signal blk00000003_sig0000009e : STD_LOGIC; 
  signal blk00000003_sig0000009d : STD_LOGIC; 
  signal blk00000003_sig0000009c : STD_LOGIC; 
  signal blk00000003_sig0000009b : STD_LOGIC; 
  signal blk00000003_sig0000009a : STD_LOGIC; 
  signal blk00000003_sig00000099 : STD_LOGIC; 
  signal blk00000003_sig00000098 : STD_LOGIC; 
  signal blk00000003_sig00000097 : STD_LOGIC; 
  signal blk00000003_sig00000096 : STD_LOGIC; 
  signal blk00000003_sig00000095 : STD_LOGIC; 
  signal blk00000003_sig00000094 : STD_LOGIC; 
  signal blk00000003_sig00000093 : STD_LOGIC; 
  signal blk00000003_sig00000092 : STD_LOGIC; 
  signal blk00000003_sig00000091 : STD_LOGIC; 
  signal blk00000003_sig00000090 : STD_LOGIC; 
  signal blk00000003_sig0000008f : STD_LOGIC; 
  signal blk00000003_sig0000008e : STD_LOGIC; 
  signal blk00000003_sig0000008d : STD_LOGIC; 
  signal blk00000003_sig0000008c : STD_LOGIC; 
  signal blk00000003_sig0000008b : STD_LOGIC; 
  signal blk00000003_sig0000008a : STD_LOGIC; 
  signal blk00000003_sig00000089 : STD_LOGIC; 
  signal blk00000003_sig00000088 : STD_LOGIC; 
  signal blk00000003_sig00000087 : STD_LOGIC; 
  signal blk00000003_sig00000086 : STD_LOGIC; 
  signal blk00000003_sig00000085 : STD_LOGIC; 
  signal blk00000003_sig00000084 : STD_LOGIC; 
  signal blk00000003_sig00000083 : STD_LOGIC; 
  signal blk00000003_sig00000082 : STD_LOGIC; 
  signal blk00000003_sig00000081 : STD_LOGIC; 
  signal blk00000003_sig00000080 : STD_LOGIC; 
  signal blk00000003_sig0000007f : STD_LOGIC; 
  signal blk00000003_sig0000007e : STD_LOGIC; 
  signal blk00000003_sig0000007d : STD_LOGIC; 
  signal blk00000003_sig0000007c : STD_LOGIC; 
  signal blk00000003_sig0000007b : STD_LOGIC; 
  signal blk00000003_sig0000007a : STD_LOGIC; 
  signal blk00000003_sig00000079 : STD_LOGIC; 
  signal blk00000003_sig00000078 : STD_LOGIC; 
  signal blk00000003_sig00000077 : STD_LOGIC; 
  signal blk00000003_sig00000076 : STD_LOGIC; 
  signal blk00000003_sig00000075 : STD_LOGIC; 
  signal blk00000003_sig00000074 : STD_LOGIC; 
  signal blk00000003_sig00000073 : STD_LOGIC; 
  signal blk00000003_sig00000072 : STD_LOGIC; 
  signal blk00000003_sig00000071 : STD_LOGIC; 
  signal blk00000003_sig00000070 : STD_LOGIC; 
  signal blk00000003_sig0000006f : STD_LOGIC; 
  signal blk00000003_sig0000006e : STD_LOGIC; 
  signal blk00000003_sig0000006d : STD_LOGIC; 
  signal blk00000003_sig0000006c : STD_LOGIC; 
  signal blk00000003_sig0000006b : STD_LOGIC; 
  signal blk00000003_sig0000006a : STD_LOGIC; 
  signal blk00000003_sig00000069 : STD_LOGIC; 
  signal blk00000003_sig00000068 : STD_LOGIC; 
  signal blk00000003_sig00000067 : STD_LOGIC; 
  signal blk00000003_sig00000066 : STD_LOGIC; 
  signal blk00000003_sig00000065 : STD_LOGIC; 
  signal blk00000003_sig00000064 : STD_LOGIC; 
  signal blk00000003_sig00000063 : STD_LOGIC; 
  signal blk00000003_sig00000062 : STD_LOGIC; 
  signal blk00000003_sig00000061 : STD_LOGIC; 
  signal blk00000003_sig00000060 : STD_LOGIC; 
  signal blk00000003_sig0000005f : STD_LOGIC; 
  signal blk00000003_sig0000005e : STD_LOGIC; 
  signal blk00000003_sig0000005d : STD_LOGIC; 
  signal blk00000003_sig0000005c : STD_LOGIC; 
  signal blk00000003_sig0000005b : STD_LOGIC; 
  signal blk00000003_sig0000005a : STD_LOGIC; 
  signal blk00000003_sig00000059 : STD_LOGIC; 
  signal blk00000003_sig00000058 : STD_LOGIC; 
  signal blk00000003_sig00000057 : STD_LOGIC; 
  signal blk00000003_sig00000056 : STD_LOGIC; 
  signal blk00000003_sig00000055 : STD_LOGIC; 
  signal blk00000003_sig00000054 : STD_LOGIC; 
  signal blk00000003_sig00000053 : STD_LOGIC; 
  signal blk00000003_sig00000052 : STD_LOGIC; 
  signal blk00000003_sig00000051 : STD_LOGIC; 
  signal blk00000003_sig00000050 : STD_LOGIC; 
  signal blk00000003_sig0000004f : STD_LOGIC; 
  signal blk00000003_sig0000004e : STD_LOGIC; 
  signal blk00000003_sig0000004d : STD_LOGIC; 
  signal blk00000003_sig0000004c : STD_LOGIC; 
  signal blk00000003_sig0000004b : STD_LOGIC; 
  signal blk00000003_sig0000004a : STD_LOGIC; 
  signal blk00000003_sig00000049 : STD_LOGIC; 
  signal blk00000003_sig00000048 : STD_LOGIC; 
  signal blk00000003_sig00000047 : STD_LOGIC; 
  signal blk00000003_sig00000046 : STD_LOGIC; 
  signal blk00000003_sig00000045 : STD_LOGIC; 
  signal blk00000003_sig00000043 : STD_LOGIC; 
  signal NLW_blk00000001_P_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000002_G_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000003_blk0000016e_O_UNCONNECTED : STD_LOGIC; 
begin
  rfd <= NlwRenamedSig_OI_rfd;
  blk00000001 : VCC
    port map (
      P => NLW_blk00000001_P_UNCONNECTED
    );
  blk00000002 : GND
    port map (
      G => NLW_blk00000002_G_UNCONNECTED
    );
  blk00000003_blk000006e8 : INV
    port map (
      I => blk00000003_sig000001b1,
      O => blk00000003_sig000001cf
    );
  blk00000003_blk000006e7 : INV
    port map (
      I => blk00000003_sig000001b2,
      O => blk00000003_sig000001d2
    );
  blk00000003_blk000006e6 : INV
    port map (
      I => blk00000003_sig000001b3,
      O => blk00000003_sig000001d5
    );
  blk00000003_blk000006e5 : INV
    port map (
      I => blk00000003_sig000001b4,
      O => blk00000003_sig000001d8
    );
  blk00000003_blk000006e4 : INV
    port map (
      I => blk00000003_sig000001b5,
      O => blk00000003_sig000001db
    );
  blk00000003_blk000006e3 : INV
    port map (
      I => blk00000003_sig000001b6,
      O => blk00000003_sig000001de
    );
  blk00000003_blk000006e2 : INV
    port map (
      I => blk00000003_sig000001b7,
      O => blk00000003_sig000001e1
    );
  blk00000003_blk000006e1 : INV
    port map (
      I => blk00000003_sig000001b8,
      O => blk00000003_sig000001e4
    );
  blk00000003_blk000006e0 : INV
    port map (
      I => blk00000003_sig000001ab,
      O => blk00000003_sig000001bd
    );
  blk00000003_blk000006df : INV
    port map (
      I => blk00000003_sig000001ac,
      O => blk00000003_sig000001c0
    );
  blk00000003_blk000006de : INV
    port map (
      I => blk00000003_sig000001ad,
      O => blk00000003_sig000001c3
    );
  blk00000003_blk000006dd : INV
    port map (
      I => blk00000003_sig000001ae,
      O => blk00000003_sig000001c6
    );
  blk00000003_blk000006dc : INV
    port map (
      I => blk00000003_sig000001af,
      O => blk00000003_sig000001c9
    );
  blk00000003_blk000006db : INV
    port map (
      I => blk00000003_sig000001b0,
      O => blk00000003_sig000001cc
    );
  blk00000003_blk000006da : INV
    port map (
      I => blk00000003_sig000001b9,
      O => blk00000003_sig000001e7
    );
  blk00000003_blk000006d9 : INV
    port map (
      I => blk00000003_sig000006b3,
      O => blk00000003_sig0000008b
    );
  blk00000003_blk000006d8 : INV
    port map (
      I => blk00000003_sig000006b4,
      O => blk00000003_sig0000008c
    );
  blk00000003_blk000006d7 : INV
    port map (
      I => blk00000003_sig000006b5,
      O => blk00000003_sig0000008d
    );
  blk00000003_blk000006d6 : INV
    port map (
      I => blk00000003_sig000006b6,
      O => blk00000003_sig0000008e
    );
  blk00000003_blk000006d5 : INV
    port map (
      I => blk00000003_sig000006b7,
      O => blk00000003_sig0000008f
    );
  blk00000003_blk000006d4 : INV
    port map (
      I => blk00000003_sig000006b8,
      O => blk00000003_sig00000090
    );
  blk00000003_blk000006d3 : INV
    port map (
      I => blk00000003_sig000006b9,
      O => blk00000003_sig00000091
    );
  blk00000003_blk000006d2 : INV
    port map (
      I => blk00000003_sig000006ba,
      O => blk00000003_sig00000092
    );
  blk00000003_blk000006d1 : INV
    port map (
      I => blk00000003_sig000006bb,
      O => blk00000003_sig00000093
    );
  blk00000003_blk000006d0 : INV
    port map (
      I => blk00000003_sig000006bc,
      O => blk00000003_sig00000094
    );
  blk00000003_blk000006cf : INV
    port map (
      I => blk00000003_sig000006bd,
      O => blk00000003_sig00000095
    );
  blk00000003_blk000006ce : INV
    port map (
      I => blk00000003_sig000006be,
      O => blk00000003_sig00000096
    );
  blk00000003_blk000006cd : INV
    port map (
      I => blk00000003_sig000006bf,
      O => blk00000003_sig00000097
    );
  blk00000003_blk000006cc : INV
    port map (
      I => blk00000003_sig000006c0,
      O => blk00000003_sig00000098
    );
  blk00000003_blk000006cb : INV
    port map (
      I => blk00000003_sig000006c1,
      O => blk00000003_sig00000099
    );
  blk00000003_blk000006ca : INV
    port map (
      I => blk00000003_sig00000611,
      O => blk00000003_sig000005fc
    );
  blk00000003_blk000006c9 : INV
    port map (
      I => blk00000003_sig00000612,
      O => blk00000003_sig000005b7
    );
  blk00000003_blk000006c8 : INV
    port map (
      I => blk00000003_sig00000613,
      O => blk00000003_sig00000572
    );
  blk00000003_blk000006c7 : INV
    port map (
      I => blk00000003_sig00000614,
      O => blk00000003_sig0000052d
    );
  blk00000003_blk000006c6 : INV
    port map (
      I => blk00000003_sig00000615,
      O => blk00000003_sig000004e8
    );
  blk00000003_blk000006c5 : INV
    port map (
      I => blk00000003_sig00000616,
      O => blk00000003_sig000004a3
    );
  blk00000003_blk000006c4 : INV
    port map (
      I => blk00000003_sig00000617,
      O => blk00000003_sig0000045e
    );
  blk00000003_blk000006c3 : INV
    port map (
      I => blk00000003_sig00000618,
      O => blk00000003_sig00000418
    );
  blk00000003_blk000006c2 : INV
    port map (
      I => blk00000003_sig00000067,
      O => blk00000003_sig000003d2
    );
  blk00000003_blk000006c1 : INV
    port map (
      I => blk00000003_sig00000075,
      O => blk00000003_sig0000038c
    );
  blk00000003_blk000006c0 : INV
    port map (
      I => blk00000003_sig0000007b,
      O => blk00000003_sig00000346
    );
  blk00000003_blk000006bf : INV
    port map (
      I => blk00000003_sig00000080,
      O => blk00000003_sig00000300
    );
  blk00000003_blk000006be : INV
    port map (
      I => blk00000003_sig00000084,
      O => blk00000003_sig000002ba
    );
  blk00000003_blk000006bd : INV
    port map (
      I => blk00000003_sig00000087,
      O => blk00000003_sig00000274
    );
  blk00000003_blk000006bc : INV
    port map (
      I => blk00000003_sig00000089,
      O => blk00000003_sig0000022e
    );
  blk00000003_blk000006bb : LUT1
    generic map(
      INIT => X"1"
    )
    port map (
      I0 => blk00000003_sig000001ec,
      O => blk00000003_sig00000089
    );
  blk00000003_blk000006ba : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000607,
      I1 => blk00000003_sig000000b8,
      I2 => blk00000003_sig00000600,
      O => blk00000003_sig000006d5
    );
  blk00000003_blk000006b9 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000608,
      I1 => blk00000003_sig000000ba,
      I2 => blk00000003_sig00000600,
      O => blk00000003_sig000006d8
    );
  blk00000003_blk000006b8 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000609,
      I1 => blk00000003_sig000000bc,
      I2 => blk00000003_sig00000600,
      O => blk00000003_sig000006db
    );
  blk00000003_blk000006b7 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig0000060a,
      I1 => blk00000003_sig000000be,
      I2 => blk00000003_sig00000600,
      O => blk00000003_sig000006de
    );
  blk00000003_blk000006b6 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig0000060b,
      I1 => blk00000003_sig000000c0,
      I2 => blk00000003_sig00000600,
      O => blk00000003_sig000006e1
    );
  blk00000003_blk000006b5 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig0000060c,
      I1 => blk00000003_sig000000c2,
      I2 => blk00000003_sig00000600,
      O => blk00000003_sig000006e4
    );
  blk00000003_blk000006b4 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig0000060d,
      I1 => blk00000003_sig000000c4,
      I2 => blk00000003_sig00000600,
      O => blk00000003_sig000006e7
    );
  blk00000003_blk000006b3 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig0000060e,
      I1 => blk00000003_sig000000c6,
      I2 => blk00000003_sig00000600,
      O => blk00000003_sig000006ea
    );
  blk00000003_blk000006b2 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000601,
      I1 => blk00000003_sig000000ac,
      I2 => blk00000003_sig00000600,
      O => blk00000003_sig000006c3
    );
  blk00000003_blk000006b1 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000602,
      I1 => blk00000003_sig000000ae,
      I2 => blk00000003_sig00000600,
      O => blk00000003_sig000006c6
    );
  blk00000003_blk000006b0 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000603,
      I1 => blk00000003_sig000000b0,
      I2 => blk00000003_sig00000600,
      O => blk00000003_sig000006c9
    );
  blk00000003_blk000006af : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000604,
      I1 => blk00000003_sig000000b2,
      I2 => blk00000003_sig00000600,
      O => blk00000003_sig000006cc
    );
  blk00000003_blk000006ae : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000605,
      I1 => blk00000003_sig000000b4,
      I2 => blk00000003_sig00000600,
      O => blk00000003_sig000006cf
    );
  blk00000003_blk000006ad : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000606,
      I1 => blk00000003_sig000000b6,
      I2 => blk00000003_sig00000600,
      O => blk00000003_sig000006d2
    );
  blk00000003_blk000006ac : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig0000060f,
      I1 => blk00000003_sig000000c8,
      I2 => blk00000003_sig00000600,
      O => blk00000003_sig000006ed
    );
  blk00000003_blk000006ab : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000610,
      I1 => blk00000003_sig000000ca,
      I2 => blk00000003_sig00000600,
      O => blk00000003_sig00000702
    );
  blk00000003_blk000006aa : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005f1,
      I1 => blk00000003_sig000000b7,
      I2 => blk00000003_sig00000611,
      O => blk00000003_sig000005d1
    );
  blk00000003_blk000006a9 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005f2,
      I1 => blk00000003_sig000000b9,
      I2 => blk00000003_sig00000611,
      O => blk00000003_sig000005d4
    );
  blk00000003_blk000006a8 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005f3,
      I1 => blk00000003_sig000000bb,
      I2 => blk00000003_sig00000611,
      O => blk00000003_sig000005d7
    );
  blk00000003_blk000006a7 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005f4,
      I1 => blk00000003_sig000000bd,
      I2 => blk00000003_sig00000611,
      O => blk00000003_sig000005da
    );
  blk00000003_blk000006a6 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005f5,
      I1 => blk00000003_sig000000bf,
      I2 => blk00000003_sig00000611,
      O => blk00000003_sig000005dd
    );
  blk00000003_blk000006a5 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005f6,
      I1 => blk00000003_sig000000c1,
      I2 => blk00000003_sig00000611,
      O => blk00000003_sig000005e0
    );
  blk00000003_blk000006a4 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005f7,
      I1 => blk00000003_sig000000c3,
      I2 => blk00000003_sig00000611,
      O => blk00000003_sig000005e3
    );
  blk00000003_blk000006a3 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005f8,
      I1 => blk00000003_sig000000c5,
      I2 => blk00000003_sig00000611,
      O => blk00000003_sig000005e6
    );
  blk00000003_blk000006a2 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000005fa,
      I1 => blk00000003_sig00000611,
      O => blk00000003_sig000005bc
    );
  blk00000003_blk000006a1 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005eb,
      I1 => blk00000003_sig000000ab,
      I2 => blk00000003_sig00000611,
      O => blk00000003_sig000005bf
    );
  blk00000003_blk000006a0 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005ec,
      I1 => blk00000003_sig000000ad,
      I2 => blk00000003_sig00000611,
      O => blk00000003_sig000005c2
    );
  blk00000003_blk0000069f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005ed,
      I1 => blk00000003_sig000000af,
      I2 => blk00000003_sig00000611,
      O => blk00000003_sig000005c5
    );
  blk00000003_blk0000069e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005ee,
      I1 => blk00000003_sig000000b1,
      I2 => blk00000003_sig00000611,
      O => blk00000003_sig000005c8
    );
  blk00000003_blk0000069d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005ef,
      I1 => blk00000003_sig000000b3,
      I2 => blk00000003_sig00000611,
      O => blk00000003_sig000005cb
    );
  blk00000003_blk0000069c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005f0,
      I1 => blk00000003_sig000000b5,
      I2 => blk00000003_sig00000611,
      O => blk00000003_sig000005ce
    );
  blk00000003_blk0000069b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005f9,
      I1 => blk00000003_sig000000c7,
      I2 => blk00000003_sig00000611,
      O => blk00000003_sig000005e9
    );
  blk00000003_blk0000069a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000008a,
      I1 => blk00000003_sig000000c9,
      I2 => blk00000003_sig00000611,
      O => blk00000003_sig000005fd
    );
  blk00000003_blk00000699 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005ac,
      I1 => blk00000003_sig000000d1,
      I2 => blk00000003_sig00000612,
      O => blk00000003_sig0000058c
    );
  blk00000003_blk00000698 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005ad,
      I1 => blk00000003_sig000000d2,
      I2 => blk00000003_sig00000612,
      O => blk00000003_sig0000058f
    );
  blk00000003_blk00000697 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005ae,
      I1 => blk00000003_sig000000d3,
      I2 => blk00000003_sig00000612,
      O => blk00000003_sig00000592
    );
  blk00000003_blk00000696 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005af,
      I1 => blk00000003_sig000000d4,
      I2 => blk00000003_sig00000612,
      O => blk00000003_sig00000595
    );
  blk00000003_blk00000695 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005b0,
      I1 => blk00000003_sig000000d5,
      I2 => blk00000003_sig00000612,
      O => blk00000003_sig00000598
    );
  blk00000003_blk00000694 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005b1,
      I1 => blk00000003_sig000000d6,
      I2 => blk00000003_sig00000612,
      O => blk00000003_sig0000059b
    );
  blk00000003_blk00000693 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005b2,
      I1 => blk00000003_sig000000d7,
      I2 => blk00000003_sig00000612,
      O => blk00000003_sig0000059e
    );
  blk00000003_blk00000692 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005b3,
      I1 => blk00000003_sig000000d8,
      I2 => blk00000003_sig00000612,
      O => blk00000003_sig000005a1
    );
  blk00000003_blk00000691 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000005b5,
      I1 => blk00000003_sig00000612,
      O => blk00000003_sig00000577
    );
  blk00000003_blk00000690 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005a6,
      I1 => blk00000003_sig000000cb,
      I2 => blk00000003_sig00000612,
      O => blk00000003_sig0000057a
    );
  blk00000003_blk0000068f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005a7,
      I1 => blk00000003_sig000000cc,
      I2 => blk00000003_sig00000612,
      O => blk00000003_sig0000057d
    );
  blk00000003_blk0000068e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005a8,
      I1 => blk00000003_sig000000cd,
      I2 => blk00000003_sig00000612,
      O => blk00000003_sig00000580
    );
  blk00000003_blk0000068d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005a9,
      I1 => blk00000003_sig000000ce,
      I2 => blk00000003_sig00000612,
      O => blk00000003_sig00000583
    );
  blk00000003_blk0000068c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005aa,
      I1 => blk00000003_sig000000cf,
      I2 => blk00000003_sig00000612,
      O => blk00000003_sig00000586
    );
  blk00000003_blk0000068b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005ab,
      I1 => blk00000003_sig000000d0,
      I2 => blk00000003_sig00000612,
      O => blk00000003_sig00000589
    );
  blk00000003_blk0000068a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005b4,
      I1 => blk00000003_sig000000d9,
      I2 => blk00000003_sig00000612,
      O => blk00000003_sig000005a4
    );
  blk00000003_blk00000689 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000048,
      I1 => blk00000003_sig000000da,
      I2 => blk00000003_sig00000612,
      O => blk00000003_sig000005b8
    );
  blk00000003_blk00000688 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000567,
      I1 => blk00000003_sig000000e1,
      I2 => blk00000003_sig00000613,
      O => blk00000003_sig00000547
    );
  blk00000003_blk00000687 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000568,
      I1 => blk00000003_sig000000e2,
      I2 => blk00000003_sig00000613,
      O => blk00000003_sig0000054a
    );
  blk00000003_blk00000686 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000569,
      I1 => blk00000003_sig000000e3,
      I2 => blk00000003_sig00000613,
      O => blk00000003_sig0000054d
    );
  blk00000003_blk00000685 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000056a,
      I1 => blk00000003_sig000000e4,
      I2 => blk00000003_sig00000613,
      O => blk00000003_sig00000550
    );
  blk00000003_blk00000684 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000056b,
      I1 => blk00000003_sig000000e5,
      I2 => blk00000003_sig00000613,
      O => blk00000003_sig00000553
    );
  blk00000003_blk00000683 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000056c,
      I1 => blk00000003_sig000000e6,
      I2 => blk00000003_sig00000613,
      O => blk00000003_sig00000556
    );
  blk00000003_blk00000682 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000056d,
      I1 => blk00000003_sig000000e7,
      I2 => blk00000003_sig00000613,
      O => blk00000003_sig00000559
    );
  blk00000003_blk00000681 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000056e,
      I1 => blk00000003_sig000000e8,
      I2 => blk00000003_sig00000613,
      O => blk00000003_sig0000055c
    );
  blk00000003_blk00000680 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000570,
      I1 => blk00000003_sig00000613,
      O => blk00000003_sig00000532
    );
  blk00000003_blk0000067f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000561,
      I1 => blk00000003_sig000000db,
      I2 => blk00000003_sig00000613,
      O => blk00000003_sig00000535
    );
  blk00000003_blk0000067e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000562,
      I1 => blk00000003_sig000000dc,
      I2 => blk00000003_sig00000613,
      O => blk00000003_sig00000538
    );
  blk00000003_blk0000067d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000563,
      I1 => blk00000003_sig000000dd,
      I2 => blk00000003_sig00000613,
      O => blk00000003_sig0000053b
    );
  blk00000003_blk0000067c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000564,
      I1 => blk00000003_sig000000de,
      I2 => blk00000003_sig00000613,
      O => blk00000003_sig0000053e
    );
  blk00000003_blk0000067b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000565,
      I1 => blk00000003_sig000000df,
      I2 => blk00000003_sig00000613,
      O => blk00000003_sig00000541
    );
  blk00000003_blk0000067a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000566,
      I1 => blk00000003_sig000000e0,
      I2 => blk00000003_sig00000613,
      O => blk00000003_sig00000544
    );
  blk00000003_blk00000679 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000056f,
      I1 => blk00000003_sig000000e9,
      I2 => blk00000003_sig00000613,
      O => blk00000003_sig0000055f
    );
  blk00000003_blk00000678 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000004c,
      I1 => blk00000003_sig000000ea,
      I2 => blk00000003_sig00000613,
      O => blk00000003_sig00000573
    );
  blk00000003_blk00000677 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000522,
      I1 => blk00000003_sig000000f1,
      I2 => blk00000003_sig00000614,
      O => blk00000003_sig00000502
    );
  blk00000003_blk00000676 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000523,
      I1 => blk00000003_sig000000f2,
      I2 => blk00000003_sig00000614,
      O => blk00000003_sig00000505
    );
  blk00000003_blk00000675 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000524,
      I1 => blk00000003_sig000000f3,
      I2 => blk00000003_sig00000614,
      O => blk00000003_sig00000508
    );
  blk00000003_blk00000674 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000525,
      I1 => blk00000003_sig000000f4,
      I2 => blk00000003_sig00000614,
      O => blk00000003_sig0000050b
    );
  blk00000003_blk00000673 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000526,
      I1 => blk00000003_sig000000f5,
      I2 => blk00000003_sig00000614,
      O => blk00000003_sig0000050e
    );
  blk00000003_blk00000672 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000527,
      I1 => blk00000003_sig000000f6,
      I2 => blk00000003_sig00000614,
      O => blk00000003_sig00000511
    );
  blk00000003_blk00000671 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000528,
      I1 => blk00000003_sig000000f7,
      I2 => blk00000003_sig00000614,
      O => blk00000003_sig00000514
    );
  blk00000003_blk00000670 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000529,
      I1 => blk00000003_sig000000f8,
      I2 => blk00000003_sig00000614,
      O => blk00000003_sig00000517
    );
  blk00000003_blk0000066f : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000052b,
      I1 => blk00000003_sig00000614,
      O => blk00000003_sig000004ed
    );
  blk00000003_blk0000066e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000051c,
      I1 => blk00000003_sig000000eb,
      I2 => blk00000003_sig00000614,
      O => blk00000003_sig000004f0
    );
  blk00000003_blk0000066d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000051d,
      I1 => blk00000003_sig000000ec,
      I2 => blk00000003_sig00000614,
      O => blk00000003_sig000004f3
    );
  blk00000003_blk0000066c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000051e,
      I1 => blk00000003_sig000000ed,
      I2 => blk00000003_sig00000614,
      O => blk00000003_sig000004f6
    );
  blk00000003_blk0000066b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000051f,
      I1 => blk00000003_sig000000ee,
      I2 => blk00000003_sig00000614,
      O => blk00000003_sig000004f9
    );
  blk00000003_blk0000066a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000520,
      I1 => blk00000003_sig000000ef,
      I2 => blk00000003_sig00000614,
      O => blk00000003_sig000004fc
    );
  blk00000003_blk00000669 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000521,
      I1 => blk00000003_sig000000f0,
      I2 => blk00000003_sig00000614,
      O => blk00000003_sig000004ff
    );
  blk00000003_blk00000668 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000052a,
      I1 => blk00000003_sig000000f9,
      I2 => blk00000003_sig00000614,
      O => blk00000003_sig0000051a
    );
  blk00000003_blk00000667 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000051,
      I1 => blk00000003_sig000000fa,
      I2 => blk00000003_sig00000614,
      O => blk00000003_sig0000052e
    );
  blk00000003_blk00000666 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004dd,
      I1 => blk00000003_sig00000101,
      I2 => blk00000003_sig00000615,
      O => blk00000003_sig000004bd
    );
  blk00000003_blk00000665 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004de,
      I1 => blk00000003_sig00000102,
      I2 => blk00000003_sig00000615,
      O => blk00000003_sig000004c0
    );
  blk00000003_blk00000664 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004df,
      I1 => blk00000003_sig00000103,
      I2 => blk00000003_sig00000615,
      O => blk00000003_sig000004c3
    );
  blk00000003_blk00000663 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004e0,
      I1 => blk00000003_sig00000104,
      I2 => blk00000003_sig00000615,
      O => blk00000003_sig000004c6
    );
  blk00000003_blk00000662 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004e1,
      I1 => blk00000003_sig00000105,
      I2 => blk00000003_sig00000615,
      O => blk00000003_sig000004c9
    );
  blk00000003_blk00000661 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004e2,
      I1 => blk00000003_sig00000106,
      I2 => blk00000003_sig00000615,
      O => blk00000003_sig000004cc
    );
  blk00000003_blk00000660 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004e3,
      I1 => blk00000003_sig00000107,
      I2 => blk00000003_sig00000615,
      O => blk00000003_sig000004cf
    );
  blk00000003_blk0000065f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004e4,
      I1 => blk00000003_sig00000108,
      I2 => blk00000003_sig00000615,
      O => blk00000003_sig000004d2
    );
  blk00000003_blk0000065e : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000004e6,
      I1 => blk00000003_sig00000615,
      O => blk00000003_sig000004a8
    );
  blk00000003_blk0000065d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004d7,
      I1 => blk00000003_sig000000fb,
      I2 => blk00000003_sig00000615,
      O => blk00000003_sig000004ab
    );
  blk00000003_blk0000065c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004d8,
      I1 => blk00000003_sig000000fc,
      I2 => blk00000003_sig00000615,
      O => blk00000003_sig000004ae
    );
  blk00000003_blk0000065b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004d9,
      I1 => blk00000003_sig000000fd,
      I2 => blk00000003_sig00000615,
      O => blk00000003_sig000004b1
    );
  blk00000003_blk0000065a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004da,
      I1 => blk00000003_sig000000fe,
      I2 => blk00000003_sig00000615,
      O => blk00000003_sig000004b4
    );
  blk00000003_blk00000659 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004db,
      I1 => blk00000003_sig000000ff,
      I2 => blk00000003_sig00000615,
      O => blk00000003_sig000004b7
    );
  blk00000003_blk00000658 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004dc,
      I1 => blk00000003_sig00000100,
      I2 => blk00000003_sig00000615,
      O => blk00000003_sig000004ba
    );
  blk00000003_blk00000657 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004e5,
      I1 => blk00000003_sig00000109,
      I2 => blk00000003_sig00000615,
      O => blk00000003_sig000004d5
    );
  blk00000003_blk00000656 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000057,
      I1 => blk00000003_sig0000010a,
      I2 => blk00000003_sig00000615,
      O => blk00000003_sig000004e9
    );
  blk00000003_blk00000655 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000498,
      I1 => blk00000003_sig00000111,
      I2 => blk00000003_sig00000616,
      O => blk00000003_sig00000478
    );
  blk00000003_blk00000654 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000499,
      I1 => blk00000003_sig00000112,
      I2 => blk00000003_sig00000616,
      O => blk00000003_sig0000047b
    );
  blk00000003_blk00000653 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000049a,
      I1 => blk00000003_sig00000113,
      I2 => blk00000003_sig00000616,
      O => blk00000003_sig0000047e
    );
  blk00000003_blk00000652 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000049b,
      I1 => blk00000003_sig00000114,
      I2 => blk00000003_sig00000616,
      O => blk00000003_sig00000481
    );
  blk00000003_blk00000651 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000049c,
      I1 => blk00000003_sig00000115,
      I2 => blk00000003_sig00000616,
      O => blk00000003_sig00000484
    );
  blk00000003_blk00000650 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000049d,
      I1 => blk00000003_sig00000116,
      I2 => blk00000003_sig00000616,
      O => blk00000003_sig00000487
    );
  blk00000003_blk0000064f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000049e,
      I1 => blk00000003_sig00000117,
      I2 => blk00000003_sig00000616,
      O => blk00000003_sig0000048a
    );
  blk00000003_blk0000064e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000049f,
      I1 => blk00000003_sig00000118,
      I2 => blk00000003_sig00000616,
      O => blk00000003_sig0000048d
    );
  blk00000003_blk0000064d : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000004a1,
      I1 => blk00000003_sig00000616,
      O => blk00000003_sig00000463
    );
  blk00000003_blk0000064c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000492,
      I1 => blk00000003_sig0000010b,
      I2 => blk00000003_sig00000616,
      O => blk00000003_sig00000466
    );
  blk00000003_blk0000064b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000493,
      I1 => blk00000003_sig0000010c,
      I2 => blk00000003_sig00000616,
      O => blk00000003_sig00000469
    );
  blk00000003_blk0000064a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000494,
      I1 => blk00000003_sig0000010d,
      I2 => blk00000003_sig00000616,
      O => blk00000003_sig0000046c
    );
  blk00000003_blk00000649 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000495,
      I1 => blk00000003_sig0000010e,
      I2 => blk00000003_sig00000616,
      O => blk00000003_sig0000046f
    );
  blk00000003_blk00000648 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000496,
      I1 => blk00000003_sig0000010f,
      I2 => blk00000003_sig00000616,
      O => blk00000003_sig00000472
    );
  blk00000003_blk00000647 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000497,
      I1 => blk00000003_sig00000110,
      I2 => blk00000003_sig00000616,
      O => blk00000003_sig00000475
    );
  blk00000003_blk00000646 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004a0,
      I1 => blk00000003_sig00000119,
      I2 => blk00000003_sig00000616,
      O => blk00000003_sig00000490
    );
  blk00000003_blk00000645 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000005e,
      I1 => blk00000003_sig0000011a,
      I2 => blk00000003_sig00000616,
      O => blk00000003_sig000004a4
    );
  blk00000003_blk00000644 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000453,
      I1 => blk00000003_sig00000121,
      I2 => blk00000003_sig00000617,
      O => blk00000003_sig00000433
    );
  blk00000003_blk00000643 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000454,
      I1 => blk00000003_sig00000122,
      I2 => blk00000003_sig00000617,
      O => blk00000003_sig00000436
    );
  blk00000003_blk00000642 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000455,
      I1 => blk00000003_sig00000123,
      I2 => blk00000003_sig00000617,
      O => blk00000003_sig00000439
    );
  blk00000003_blk00000641 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000456,
      I1 => blk00000003_sig00000124,
      I2 => blk00000003_sig00000617,
      O => blk00000003_sig0000043c
    );
  blk00000003_blk00000640 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000457,
      I1 => blk00000003_sig00000125,
      I2 => blk00000003_sig00000617,
      O => blk00000003_sig0000043f
    );
  blk00000003_blk0000063f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000458,
      I1 => blk00000003_sig00000126,
      I2 => blk00000003_sig00000617,
      O => blk00000003_sig00000442
    );
  blk00000003_blk0000063e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000459,
      I1 => blk00000003_sig00000127,
      I2 => blk00000003_sig00000617,
      O => blk00000003_sig00000445
    );
  blk00000003_blk0000063d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000045a,
      I1 => blk00000003_sig00000128,
      I2 => blk00000003_sig00000617,
      O => blk00000003_sig00000448
    );
  blk00000003_blk0000063c : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000045c,
      I1 => blk00000003_sig00000617,
      O => blk00000003_sig0000041e
    );
  blk00000003_blk0000063b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000044d,
      I1 => blk00000003_sig0000011b,
      I2 => blk00000003_sig00000617,
      O => blk00000003_sig00000421
    );
  blk00000003_blk0000063a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000044e,
      I1 => blk00000003_sig0000011c,
      I2 => blk00000003_sig00000617,
      O => blk00000003_sig00000424
    );
  blk00000003_blk00000639 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000044f,
      I1 => blk00000003_sig0000011d,
      I2 => blk00000003_sig00000617,
      O => blk00000003_sig00000427
    );
  blk00000003_blk00000638 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000450,
      I1 => blk00000003_sig0000011e,
      I2 => blk00000003_sig00000617,
      O => blk00000003_sig0000042a
    );
  blk00000003_blk00000637 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000451,
      I1 => blk00000003_sig0000011f,
      I2 => blk00000003_sig00000617,
      O => blk00000003_sig0000042d
    );
  blk00000003_blk00000636 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000452,
      I1 => blk00000003_sig00000120,
      I2 => blk00000003_sig00000617,
      O => blk00000003_sig00000430
    );
  blk00000003_blk00000635 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000045b,
      I1 => blk00000003_sig00000129,
      I2 => blk00000003_sig00000617,
      O => blk00000003_sig0000044b
    );
  blk00000003_blk00000634 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000066,
      I1 => blk00000003_sig0000012a,
      I2 => blk00000003_sig00000617,
      O => blk00000003_sig0000045f
    );
  blk00000003_blk00000633 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000040d,
      I1 => blk00000003_sig00000131,
      I2 => blk00000003_sig00000618,
      O => blk00000003_sig000003ed
    );
  blk00000003_blk00000632 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000040e,
      I1 => blk00000003_sig00000132,
      I2 => blk00000003_sig00000618,
      O => blk00000003_sig000003f0
    );
  blk00000003_blk00000631 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000040f,
      I1 => blk00000003_sig00000133,
      I2 => blk00000003_sig00000618,
      O => blk00000003_sig000003f3
    );
  blk00000003_blk00000630 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000410,
      I1 => blk00000003_sig00000134,
      I2 => blk00000003_sig00000618,
      O => blk00000003_sig000003f6
    );
  blk00000003_blk0000062f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000411,
      I1 => blk00000003_sig00000135,
      I2 => blk00000003_sig00000618,
      O => blk00000003_sig000003f9
    );
  blk00000003_blk0000062e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000412,
      I1 => blk00000003_sig00000136,
      I2 => blk00000003_sig00000618,
      O => blk00000003_sig000003fc
    );
  blk00000003_blk0000062d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000413,
      I1 => blk00000003_sig00000137,
      I2 => blk00000003_sig00000618,
      O => blk00000003_sig000003ff
    );
  blk00000003_blk0000062c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000414,
      I1 => blk00000003_sig00000138,
      I2 => blk00000003_sig00000618,
      O => blk00000003_sig00000402
    );
  blk00000003_blk0000062b : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000416,
      I1 => blk00000003_sig00000618,
      O => blk00000003_sig000003d8
    );
  blk00000003_blk0000062a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000407,
      I1 => blk00000003_sig0000012b,
      I2 => blk00000003_sig00000618,
      O => blk00000003_sig000003db
    );
  blk00000003_blk00000629 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000408,
      I1 => blk00000003_sig0000012c,
      I2 => blk00000003_sig00000618,
      O => blk00000003_sig000003de
    );
  blk00000003_blk00000628 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000409,
      I1 => blk00000003_sig0000012d,
      I2 => blk00000003_sig00000618,
      O => blk00000003_sig000003e1
    );
  blk00000003_blk00000627 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000040a,
      I1 => blk00000003_sig0000012e,
      I2 => blk00000003_sig00000618,
      O => blk00000003_sig000003e4
    );
  blk00000003_blk00000626 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000040b,
      I1 => blk00000003_sig0000012f,
      I2 => blk00000003_sig00000618,
      O => blk00000003_sig000003e7
    );
  blk00000003_blk00000625 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000040c,
      I1 => blk00000003_sig00000130,
      I2 => blk00000003_sig00000618,
      O => blk00000003_sig000003ea
    );
  blk00000003_blk00000624 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000415,
      I1 => blk00000003_sig00000139,
      I2 => blk00000003_sig00000618,
      O => blk00000003_sig00000405
    );
  blk00000003_blk00000623 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000041b,
      I1 => blk00000003_sig0000013a,
      I2 => blk00000003_sig00000618,
      O => blk00000003_sig00000419
    );
  blk00000003_blk00000622 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003c7,
      I1 => blk00000003_sig00000141,
      I2 => blk00000003_sig00000067,
      O => blk00000003_sig000003a7
    );
  blk00000003_blk00000621 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003c8,
      I1 => blk00000003_sig00000142,
      I2 => blk00000003_sig00000067,
      O => blk00000003_sig000003aa
    );
  blk00000003_blk00000620 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003c9,
      I1 => blk00000003_sig00000143,
      I2 => blk00000003_sig00000067,
      O => blk00000003_sig000003ad
    );
  blk00000003_blk0000061f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003ca,
      I1 => blk00000003_sig00000144,
      I2 => blk00000003_sig00000067,
      O => blk00000003_sig000003b0
    );
  blk00000003_blk0000061e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003cb,
      I1 => blk00000003_sig00000145,
      I2 => blk00000003_sig00000067,
      O => blk00000003_sig000003b3
    );
  blk00000003_blk0000061d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003cc,
      I1 => blk00000003_sig00000146,
      I2 => blk00000003_sig00000067,
      O => blk00000003_sig000003b6
    );
  blk00000003_blk0000061c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003cd,
      I1 => blk00000003_sig00000147,
      I2 => blk00000003_sig00000067,
      O => blk00000003_sig000003b9
    );
  blk00000003_blk0000061b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003ce,
      I1 => blk00000003_sig00000148,
      I2 => blk00000003_sig00000067,
      O => blk00000003_sig000003bc
    );
  blk00000003_blk0000061a : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000003d0,
      I1 => blk00000003_sig00000067,
      O => blk00000003_sig00000392
    );
  blk00000003_blk00000619 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003c1,
      I1 => blk00000003_sig0000013b,
      I2 => blk00000003_sig00000067,
      O => blk00000003_sig00000395
    );
  blk00000003_blk00000618 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003c2,
      I1 => blk00000003_sig0000013c,
      I2 => blk00000003_sig00000067,
      O => blk00000003_sig00000398
    );
  blk00000003_blk00000617 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003c3,
      I1 => blk00000003_sig0000013d,
      I2 => blk00000003_sig00000067,
      O => blk00000003_sig0000039b
    );
  blk00000003_blk00000616 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003c4,
      I1 => blk00000003_sig0000013e,
      I2 => blk00000003_sig00000067,
      O => blk00000003_sig0000039e
    );
  blk00000003_blk00000615 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003c5,
      I1 => blk00000003_sig0000013f,
      I2 => blk00000003_sig00000067,
      O => blk00000003_sig000003a1
    );
  blk00000003_blk00000614 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003c6,
      I1 => blk00000003_sig00000140,
      I2 => blk00000003_sig00000067,
      O => blk00000003_sig000003a4
    );
  blk00000003_blk00000613 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003cf,
      I1 => blk00000003_sig00000149,
      I2 => blk00000003_sig00000067,
      O => blk00000003_sig000003bf
    );
  blk00000003_blk00000612 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003d5,
      I1 => blk00000003_sig0000014a,
      I2 => blk00000003_sig00000067,
      O => blk00000003_sig000003d3
    );
  blk00000003_blk00000611 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000381,
      I1 => blk00000003_sig00000151,
      I2 => blk00000003_sig00000075,
      O => blk00000003_sig00000361
    );
  blk00000003_blk00000610 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000382,
      I1 => blk00000003_sig00000152,
      I2 => blk00000003_sig00000075,
      O => blk00000003_sig00000364
    );
  blk00000003_blk0000060f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000383,
      I1 => blk00000003_sig00000153,
      I2 => blk00000003_sig00000075,
      O => blk00000003_sig00000367
    );
  blk00000003_blk0000060e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000384,
      I1 => blk00000003_sig00000154,
      I2 => blk00000003_sig00000075,
      O => blk00000003_sig0000036a
    );
  blk00000003_blk0000060d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000385,
      I1 => blk00000003_sig00000155,
      I2 => blk00000003_sig00000075,
      O => blk00000003_sig0000036d
    );
  blk00000003_blk0000060c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000386,
      I1 => blk00000003_sig00000156,
      I2 => blk00000003_sig00000075,
      O => blk00000003_sig00000370
    );
  blk00000003_blk0000060b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000387,
      I1 => blk00000003_sig00000157,
      I2 => blk00000003_sig00000075,
      O => blk00000003_sig00000373
    );
  blk00000003_blk0000060a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000388,
      I1 => blk00000003_sig00000158,
      I2 => blk00000003_sig00000075,
      O => blk00000003_sig00000376
    );
  blk00000003_blk00000609 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000038a,
      I1 => blk00000003_sig00000075,
      O => blk00000003_sig0000034c
    );
  blk00000003_blk00000608 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000037b,
      I1 => blk00000003_sig0000014b,
      I2 => blk00000003_sig00000075,
      O => blk00000003_sig0000034f
    );
  blk00000003_blk00000607 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000037c,
      I1 => blk00000003_sig0000014c,
      I2 => blk00000003_sig00000075,
      O => blk00000003_sig00000352
    );
  blk00000003_blk00000606 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000037d,
      I1 => blk00000003_sig0000014d,
      I2 => blk00000003_sig00000075,
      O => blk00000003_sig00000355
    );
  blk00000003_blk00000605 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000037e,
      I1 => blk00000003_sig0000014e,
      I2 => blk00000003_sig00000075,
      O => blk00000003_sig00000358
    );
  blk00000003_blk00000604 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000037f,
      I1 => blk00000003_sig0000014f,
      I2 => blk00000003_sig00000075,
      O => blk00000003_sig0000035b
    );
  blk00000003_blk00000603 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000380,
      I1 => blk00000003_sig00000150,
      I2 => blk00000003_sig00000075,
      O => blk00000003_sig0000035e
    );
  blk00000003_blk00000602 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000389,
      I1 => blk00000003_sig00000159,
      I2 => blk00000003_sig00000075,
      O => blk00000003_sig00000379
    );
  blk00000003_blk00000601 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000038f,
      I1 => blk00000003_sig0000015a,
      I2 => blk00000003_sig00000075,
      O => blk00000003_sig0000038d
    );
  blk00000003_blk00000600 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000033b,
      I1 => blk00000003_sig00000161,
      I2 => blk00000003_sig0000007b,
      O => blk00000003_sig0000031b
    );
  blk00000003_blk000005ff : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000033c,
      I1 => blk00000003_sig00000162,
      I2 => blk00000003_sig0000007b,
      O => blk00000003_sig0000031e
    );
  blk00000003_blk000005fe : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000033d,
      I1 => blk00000003_sig00000163,
      I2 => blk00000003_sig0000007b,
      O => blk00000003_sig00000321
    );
  blk00000003_blk000005fd : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000033e,
      I1 => blk00000003_sig00000164,
      I2 => blk00000003_sig0000007b,
      O => blk00000003_sig00000324
    );
  blk00000003_blk000005fc : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000033f,
      I1 => blk00000003_sig00000165,
      I2 => blk00000003_sig0000007b,
      O => blk00000003_sig00000327
    );
  blk00000003_blk000005fb : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000340,
      I1 => blk00000003_sig00000166,
      I2 => blk00000003_sig0000007b,
      O => blk00000003_sig0000032a
    );
  blk00000003_blk000005fa : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000341,
      I1 => blk00000003_sig00000167,
      I2 => blk00000003_sig0000007b,
      O => blk00000003_sig0000032d
    );
  blk00000003_blk000005f9 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000342,
      I1 => blk00000003_sig00000168,
      I2 => blk00000003_sig0000007b,
      O => blk00000003_sig00000330
    );
  blk00000003_blk000005f8 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000344,
      I1 => blk00000003_sig0000007b,
      O => blk00000003_sig00000306
    );
  blk00000003_blk000005f7 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000335,
      I1 => blk00000003_sig0000015b,
      I2 => blk00000003_sig0000007b,
      O => blk00000003_sig00000309
    );
  blk00000003_blk000005f6 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000336,
      I1 => blk00000003_sig0000015c,
      I2 => blk00000003_sig0000007b,
      O => blk00000003_sig0000030c
    );
  blk00000003_blk000005f5 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000337,
      I1 => blk00000003_sig0000015d,
      I2 => blk00000003_sig0000007b,
      O => blk00000003_sig0000030f
    );
  blk00000003_blk000005f4 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000338,
      I1 => blk00000003_sig0000015e,
      I2 => blk00000003_sig0000007b,
      O => blk00000003_sig00000312
    );
  blk00000003_blk000005f3 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000339,
      I1 => blk00000003_sig0000015f,
      I2 => blk00000003_sig0000007b,
      O => blk00000003_sig00000315
    );
  blk00000003_blk000005f2 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000033a,
      I1 => blk00000003_sig00000160,
      I2 => blk00000003_sig0000007b,
      O => blk00000003_sig00000318
    );
  blk00000003_blk000005f1 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000343,
      I1 => blk00000003_sig00000169,
      I2 => blk00000003_sig0000007b,
      O => blk00000003_sig00000333
    );
  blk00000003_blk000005f0 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000349,
      I1 => blk00000003_sig0000016a,
      I2 => blk00000003_sig0000007b,
      O => blk00000003_sig00000347
    );
  blk00000003_blk000005ef : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002f5,
      I1 => blk00000003_sig00000171,
      I2 => blk00000003_sig00000080,
      O => blk00000003_sig000002d5
    );
  blk00000003_blk000005ee : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002f6,
      I1 => blk00000003_sig00000172,
      I2 => blk00000003_sig00000080,
      O => blk00000003_sig000002d8
    );
  blk00000003_blk000005ed : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002f7,
      I1 => blk00000003_sig00000173,
      I2 => blk00000003_sig00000080,
      O => blk00000003_sig000002db
    );
  blk00000003_blk000005ec : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002f8,
      I1 => blk00000003_sig00000174,
      I2 => blk00000003_sig00000080,
      O => blk00000003_sig000002de
    );
  blk00000003_blk000005eb : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002f9,
      I1 => blk00000003_sig00000175,
      I2 => blk00000003_sig00000080,
      O => blk00000003_sig000002e1
    );
  blk00000003_blk000005ea : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002fa,
      I1 => blk00000003_sig00000176,
      I2 => blk00000003_sig00000080,
      O => blk00000003_sig000002e4
    );
  blk00000003_blk000005e9 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002fb,
      I1 => blk00000003_sig00000177,
      I2 => blk00000003_sig00000080,
      O => blk00000003_sig000002e7
    );
  blk00000003_blk000005e8 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002fc,
      I1 => blk00000003_sig00000178,
      I2 => blk00000003_sig00000080,
      O => blk00000003_sig000002ea
    );
  blk00000003_blk000005e7 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000002fe,
      I1 => blk00000003_sig00000080,
      O => blk00000003_sig000002c0
    );
  blk00000003_blk000005e6 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002ef,
      I1 => blk00000003_sig0000016b,
      I2 => blk00000003_sig00000080,
      O => blk00000003_sig000002c3
    );
  blk00000003_blk000005e5 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002f0,
      I1 => blk00000003_sig0000016c,
      I2 => blk00000003_sig00000080,
      O => blk00000003_sig000002c6
    );
  blk00000003_blk000005e4 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002f1,
      I1 => blk00000003_sig0000016d,
      I2 => blk00000003_sig00000080,
      O => blk00000003_sig000002c9
    );
  blk00000003_blk000005e3 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002f2,
      I1 => blk00000003_sig0000016e,
      I2 => blk00000003_sig00000080,
      O => blk00000003_sig000002cc
    );
  blk00000003_blk000005e2 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002f3,
      I1 => blk00000003_sig0000016f,
      I2 => blk00000003_sig00000080,
      O => blk00000003_sig000002cf
    );
  blk00000003_blk000005e1 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002f4,
      I1 => blk00000003_sig00000170,
      I2 => blk00000003_sig00000080,
      O => blk00000003_sig000002d2
    );
  blk00000003_blk000005e0 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002fd,
      I1 => blk00000003_sig00000179,
      I2 => blk00000003_sig00000080,
      O => blk00000003_sig000002ed
    );
  blk00000003_blk000005df : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000303,
      I1 => blk00000003_sig0000017a,
      I2 => blk00000003_sig00000080,
      O => blk00000003_sig00000301
    );
  blk00000003_blk000005de : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002af,
      I1 => blk00000003_sig00000181,
      I2 => blk00000003_sig00000084,
      O => blk00000003_sig0000028f
    );
  blk00000003_blk000005dd : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002b0,
      I1 => blk00000003_sig00000182,
      I2 => blk00000003_sig00000084,
      O => blk00000003_sig00000292
    );
  blk00000003_blk000005dc : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002b1,
      I1 => blk00000003_sig00000183,
      I2 => blk00000003_sig00000084,
      O => blk00000003_sig00000295
    );
  blk00000003_blk000005db : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002b2,
      I1 => blk00000003_sig00000184,
      I2 => blk00000003_sig00000084,
      O => blk00000003_sig00000298
    );
  blk00000003_blk000005da : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002b3,
      I1 => blk00000003_sig00000185,
      I2 => blk00000003_sig00000084,
      O => blk00000003_sig0000029b
    );
  blk00000003_blk000005d9 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002b4,
      I1 => blk00000003_sig00000186,
      I2 => blk00000003_sig00000084,
      O => blk00000003_sig0000029e
    );
  blk00000003_blk000005d8 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002b5,
      I1 => blk00000003_sig00000187,
      I2 => blk00000003_sig00000084,
      O => blk00000003_sig000002a1
    );
  blk00000003_blk000005d7 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002b6,
      I1 => blk00000003_sig00000188,
      I2 => blk00000003_sig00000084,
      O => blk00000003_sig000002a4
    );
  blk00000003_blk000005d6 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000002b8,
      I1 => blk00000003_sig00000084,
      O => blk00000003_sig0000027a
    );
  blk00000003_blk000005d5 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002a9,
      I1 => blk00000003_sig0000017b,
      I2 => blk00000003_sig00000084,
      O => blk00000003_sig0000027d
    );
  blk00000003_blk000005d4 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002aa,
      I1 => blk00000003_sig0000017c,
      I2 => blk00000003_sig00000084,
      O => blk00000003_sig00000280
    );
  blk00000003_blk000005d3 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002ab,
      I1 => blk00000003_sig0000017d,
      I2 => blk00000003_sig00000084,
      O => blk00000003_sig00000283
    );
  blk00000003_blk000005d2 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002ac,
      I1 => blk00000003_sig0000017e,
      I2 => blk00000003_sig00000084,
      O => blk00000003_sig00000286
    );
  blk00000003_blk000005d1 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002ad,
      I1 => blk00000003_sig0000017f,
      I2 => blk00000003_sig00000084,
      O => blk00000003_sig00000289
    );
  blk00000003_blk000005d0 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002ae,
      I1 => blk00000003_sig00000180,
      I2 => blk00000003_sig00000084,
      O => blk00000003_sig0000028c
    );
  blk00000003_blk000005cf : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002b7,
      I1 => blk00000003_sig00000189,
      I2 => blk00000003_sig00000084,
      O => blk00000003_sig000002a7
    );
  blk00000003_blk000005ce : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002bd,
      I1 => blk00000003_sig0000018a,
      I2 => blk00000003_sig00000084,
      O => blk00000003_sig000002bb
    );
  blk00000003_blk000005cd : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000269,
      I1 => blk00000003_sig00000191,
      I2 => blk00000003_sig00000087,
      O => blk00000003_sig00000249
    );
  blk00000003_blk000005cc : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000026a,
      I1 => blk00000003_sig00000192,
      I2 => blk00000003_sig00000087,
      O => blk00000003_sig0000024c
    );
  blk00000003_blk000005cb : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000026b,
      I1 => blk00000003_sig00000193,
      I2 => blk00000003_sig00000087,
      O => blk00000003_sig0000024f
    );
  blk00000003_blk000005ca : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000026c,
      I1 => blk00000003_sig00000194,
      I2 => blk00000003_sig00000087,
      O => blk00000003_sig00000252
    );
  blk00000003_blk000005c9 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000026d,
      I1 => blk00000003_sig00000195,
      I2 => blk00000003_sig00000087,
      O => blk00000003_sig00000255
    );
  blk00000003_blk000005c8 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000026e,
      I1 => blk00000003_sig00000196,
      I2 => blk00000003_sig00000087,
      O => blk00000003_sig00000258
    );
  blk00000003_blk000005c7 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000026f,
      I1 => blk00000003_sig00000197,
      I2 => blk00000003_sig00000087,
      O => blk00000003_sig0000025b
    );
  blk00000003_blk000005c6 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000270,
      I1 => blk00000003_sig00000198,
      I2 => blk00000003_sig00000087,
      O => blk00000003_sig0000025e
    );
  blk00000003_blk000005c5 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000272,
      I1 => blk00000003_sig00000087,
      O => blk00000003_sig00000234
    );
  blk00000003_blk000005c4 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000263,
      I1 => blk00000003_sig0000018b,
      I2 => blk00000003_sig00000087,
      O => blk00000003_sig00000237
    );
  blk00000003_blk000005c3 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000264,
      I1 => blk00000003_sig0000018c,
      I2 => blk00000003_sig00000087,
      O => blk00000003_sig0000023a
    );
  blk00000003_blk000005c2 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000265,
      I1 => blk00000003_sig0000018d,
      I2 => blk00000003_sig00000087,
      O => blk00000003_sig0000023d
    );
  blk00000003_blk000005c1 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000266,
      I1 => blk00000003_sig0000018e,
      I2 => blk00000003_sig00000087,
      O => blk00000003_sig00000240
    );
  blk00000003_blk000005c0 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000267,
      I1 => blk00000003_sig0000018f,
      I2 => blk00000003_sig00000087,
      O => blk00000003_sig00000243
    );
  blk00000003_blk000005bf : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000268,
      I1 => blk00000003_sig00000190,
      I2 => blk00000003_sig00000087,
      O => blk00000003_sig00000246
    );
  blk00000003_blk000005be : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000271,
      I1 => blk00000003_sig00000199,
      I2 => blk00000003_sig00000087,
      O => blk00000003_sig00000261
    );
  blk00000003_blk000005bd : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000277,
      I1 => blk00000003_sig0000019a,
      I2 => blk00000003_sig00000087,
      O => blk00000003_sig00000275
    );
  blk00000003_blk000005bc : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000223,
      I1 => blk00000003_sig000001a1,
      I2 => blk00000003_sig00000089,
      O => blk00000003_sig00000203
    );
  blk00000003_blk000005bb : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000224,
      I1 => blk00000003_sig000001a2,
      I2 => blk00000003_sig00000089,
      O => blk00000003_sig00000206
    );
  blk00000003_blk000005ba : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000225,
      I1 => blk00000003_sig000001a3,
      I2 => blk00000003_sig00000089,
      O => blk00000003_sig00000209
    );
  blk00000003_blk000005b9 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000226,
      I1 => blk00000003_sig000001a4,
      I2 => blk00000003_sig00000089,
      O => blk00000003_sig0000020c
    );
  blk00000003_blk000005b8 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000227,
      I1 => blk00000003_sig000001a5,
      I2 => blk00000003_sig00000089,
      O => blk00000003_sig0000020f
    );
  blk00000003_blk000005b7 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000228,
      I1 => blk00000003_sig000001a6,
      I2 => blk00000003_sig00000089,
      O => blk00000003_sig00000212
    );
  blk00000003_blk000005b6 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000229,
      I1 => blk00000003_sig000001a7,
      I2 => blk00000003_sig00000089,
      O => blk00000003_sig00000215
    );
  blk00000003_blk000005b5 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000022a,
      I1 => blk00000003_sig000001a8,
      I2 => blk00000003_sig00000089,
      O => blk00000003_sig00000218
    );
  blk00000003_blk000005b4 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000022c,
      I1 => blk00000003_sig00000089,
      O => blk00000003_sig000001ee
    );
  blk00000003_blk000005b3 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000021d,
      I1 => blk00000003_sig0000019b,
      I2 => blk00000003_sig00000089,
      O => blk00000003_sig000001f1
    );
  blk00000003_blk000005b2 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000021e,
      I1 => blk00000003_sig0000019c,
      I2 => blk00000003_sig00000089,
      O => blk00000003_sig000001f4
    );
  blk00000003_blk000005b1 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000021f,
      I1 => blk00000003_sig0000019d,
      I2 => blk00000003_sig00000089,
      O => blk00000003_sig000001f7
    );
  blk00000003_blk000005b0 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000220,
      I1 => blk00000003_sig0000019e,
      I2 => blk00000003_sig00000089,
      O => blk00000003_sig000001fa
    );
  blk00000003_blk000005af : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000221,
      I1 => blk00000003_sig0000019f,
      I2 => blk00000003_sig00000089,
      O => blk00000003_sig000001fd
    );
  blk00000003_blk000005ae : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000222,
      I1 => blk00000003_sig000001a0,
      I2 => blk00000003_sig00000089,
      O => blk00000003_sig00000200
    );
  blk00000003_blk000005ad : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000022b,
      I1 => blk00000003_sig000001a9,
      I2 => blk00000003_sig00000089,
      O => blk00000003_sig0000021b
    );
  blk00000003_blk000005ac : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000231,
      I1 => blk00000003_sig000001aa,
      I2 => blk00000003_sig00000089,
      O => blk00000003_sig0000022f
    );
  blk00000003_blk000005ab : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000009b,
      I1 => blk00000003_sig000001ba,
      O => blk00000003_sig000001ea
    );
  blk00000003_blk000005aa : LUT1
    generic map(
      INIT => X"1"
    )
    port map (
      I0 => blk00000003_sig00000600,
      O => blk00000003_sig0000009a
    );
  blk00000003_blk000005a9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000703,
      Q => fractional(0)
    );
  blk00000003_blk000005a8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ee,
      Q => fractional(1)
    );
  blk00000003_blk000005a7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006eb,
      Q => fractional(2)
    );
  blk00000003_blk000005a6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006e8,
      Q => fractional(3)
    );
  blk00000003_blk000005a5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006e5,
      Q => fractional(4)
    );
  blk00000003_blk000005a4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006e2,
      Q => fractional(5)
    );
  blk00000003_blk000005a3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006df,
      Q => fractional(6)
    );
  blk00000003_blk000005a2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006dc,
      Q => fractional(7)
    );
  blk00000003_blk000005a1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006d9,
      Q => fractional(8)
    );
  blk00000003_blk000005a0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006d6,
      Q => fractional(9)
    );
  blk00000003_blk0000059f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006d3,
      Q => fractional(10)
    );
  blk00000003_blk0000059e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006d0,
      Q => fractional(11)
    );
  blk00000003_blk0000059d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006cd,
      Q => fractional(12)
    );
  blk00000003_blk0000059c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ca,
      Q => fractional(13)
    );
  blk00000003_blk0000059b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006c7,
      Q => fractional(14)
    );
  blk00000003_blk0000059a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006c4,
      Q => fractional(15)
    );
  blk00000003_blk00000599 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006f0,
      Q => blk00000003_sig00000706
    );
  blk00000003_blk00000598 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006f2,
      Q => blk00000003_sig00000705
    );
  blk00000003_blk00000597 : MULT_AND
    port map (
      I0 => blk00000003_sig000000ca,
      I1 => blk00000003_sig00000600,
      LO => blk00000003_sig00000704
    );
  blk00000003_blk00000596 : MULT_AND
    port map (
      I0 => blk00000003_sig000000c8,
      I1 => blk00000003_sig00000600,
      LO => blk00000003_sig00000701
    );
  blk00000003_blk00000595 : MULT_AND
    port map (
      I0 => blk00000003_sig000000c6,
      I1 => blk00000003_sig00000600,
      LO => blk00000003_sig00000700
    );
  blk00000003_blk00000594 : MULT_AND
    port map (
      I0 => blk00000003_sig000000c4,
      I1 => blk00000003_sig00000600,
      LO => blk00000003_sig000006ff
    );
  blk00000003_blk00000593 : MULT_AND
    port map (
      I0 => blk00000003_sig000000c2,
      I1 => blk00000003_sig00000600,
      LO => blk00000003_sig000006fe
    );
  blk00000003_blk00000592 : MULT_AND
    port map (
      I0 => blk00000003_sig000000c0,
      I1 => blk00000003_sig00000600,
      LO => blk00000003_sig000006fd
    );
  blk00000003_blk00000591 : MULT_AND
    port map (
      I0 => blk00000003_sig000000be,
      I1 => blk00000003_sig00000600,
      LO => blk00000003_sig000006fc
    );
  blk00000003_blk00000590 : MULT_AND
    port map (
      I0 => blk00000003_sig000000bc,
      I1 => blk00000003_sig00000600,
      LO => blk00000003_sig000006fb
    );
  blk00000003_blk0000058f : MULT_AND
    port map (
      I0 => blk00000003_sig000000ba,
      I1 => blk00000003_sig00000600,
      LO => blk00000003_sig000006fa
    );
  blk00000003_blk0000058e : MULT_AND
    port map (
      I0 => blk00000003_sig000000b8,
      I1 => blk00000003_sig00000600,
      LO => blk00000003_sig000006f9
    );
  blk00000003_blk0000058d : MULT_AND
    port map (
      I0 => blk00000003_sig000000b6,
      I1 => blk00000003_sig00000600,
      LO => blk00000003_sig000006f8
    );
  blk00000003_blk0000058c : MULT_AND
    port map (
      I0 => blk00000003_sig000000b4,
      I1 => blk00000003_sig00000600,
      LO => blk00000003_sig000006f7
    );
  blk00000003_blk0000058b : MULT_AND
    port map (
      I0 => blk00000003_sig000000b2,
      I1 => blk00000003_sig00000600,
      LO => blk00000003_sig000006f6
    );
  blk00000003_blk0000058a : MULT_AND
    port map (
      I0 => blk00000003_sig000000b0,
      I1 => blk00000003_sig00000600,
      LO => blk00000003_sig000006f5
    );
  blk00000003_blk00000589 : MULT_AND
    port map (
      I0 => blk00000003_sig000000ae,
      I1 => blk00000003_sig00000600,
      LO => blk00000003_sig000006f4
    );
  blk00000003_blk00000588 : MULT_AND
    port map (
      I0 => blk00000003_sig000000ac,
      I1 => blk00000003_sig00000600,
      LO => blk00000003_sig000006f3
    );
  blk00000003_blk00000587 : MULT_AND
    port map (
      I0 => blk00000003_sig00000043,
      I1 => blk00000003_sig00000600,
      LO => blk00000003_sig000006f1
    );
  blk00000003_blk00000586 : MUXCY
    port map (
      CI => blk00000003_sig00000043,
      DI => blk00000003_sig00000704,
      S => blk00000003_sig00000702,
      O => blk00000003_sig000006ec
    );
  blk00000003_blk00000585 : XORCY
    port map (
      CI => blk00000003_sig00000043,
      LI => blk00000003_sig00000702,
      O => blk00000003_sig00000703
    );
  blk00000003_blk00000584 : MUXCY
    port map (
      CI => blk00000003_sig000006ec,
      DI => blk00000003_sig00000701,
      S => blk00000003_sig000006ed,
      O => blk00000003_sig000006e9
    );
  blk00000003_blk00000583 : MUXCY
    port map (
      CI => blk00000003_sig000006e9,
      DI => blk00000003_sig00000700,
      S => blk00000003_sig000006ea,
      O => blk00000003_sig000006e6
    );
  blk00000003_blk00000582 : MUXCY
    port map (
      CI => blk00000003_sig000006e6,
      DI => blk00000003_sig000006ff,
      S => blk00000003_sig000006e7,
      O => blk00000003_sig000006e3
    );
  blk00000003_blk00000581 : MUXCY
    port map (
      CI => blk00000003_sig000006e3,
      DI => blk00000003_sig000006fe,
      S => blk00000003_sig000006e4,
      O => blk00000003_sig000006e0
    );
  blk00000003_blk00000580 : MUXCY
    port map (
      CI => blk00000003_sig000006e0,
      DI => blk00000003_sig000006fd,
      S => blk00000003_sig000006e1,
      O => blk00000003_sig000006dd
    );
  blk00000003_blk0000057f : MUXCY
    port map (
      CI => blk00000003_sig000006dd,
      DI => blk00000003_sig000006fc,
      S => blk00000003_sig000006de,
      O => blk00000003_sig000006da
    );
  blk00000003_blk0000057e : MUXCY
    port map (
      CI => blk00000003_sig000006da,
      DI => blk00000003_sig000006fb,
      S => blk00000003_sig000006db,
      O => blk00000003_sig000006d7
    );
  blk00000003_blk0000057d : MUXCY
    port map (
      CI => blk00000003_sig000006d7,
      DI => blk00000003_sig000006fa,
      S => blk00000003_sig000006d8,
      O => blk00000003_sig000006d4
    );
  blk00000003_blk0000057c : MUXCY
    port map (
      CI => blk00000003_sig000006d4,
      DI => blk00000003_sig000006f9,
      S => blk00000003_sig000006d5,
      O => blk00000003_sig000006d1
    );
  blk00000003_blk0000057b : MUXCY
    port map (
      CI => blk00000003_sig000006d1,
      DI => blk00000003_sig000006f8,
      S => blk00000003_sig000006d2,
      O => blk00000003_sig000006ce
    );
  blk00000003_blk0000057a : MUXCY
    port map (
      CI => blk00000003_sig000006ce,
      DI => blk00000003_sig000006f7,
      S => blk00000003_sig000006cf,
      O => blk00000003_sig000006cb
    );
  blk00000003_blk00000579 : MUXCY
    port map (
      CI => blk00000003_sig000006cb,
      DI => blk00000003_sig000006f6,
      S => blk00000003_sig000006cc,
      O => blk00000003_sig000006c8
    );
  blk00000003_blk00000578 : MUXCY
    port map (
      CI => blk00000003_sig000006c8,
      DI => blk00000003_sig000006f5,
      S => blk00000003_sig000006c9,
      O => blk00000003_sig000006c5
    );
  blk00000003_blk00000577 : MUXCY
    port map (
      CI => blk00000003_sig000006c5,
      DI => blk00000003_sig000006f4,
      S => blk00000003_sig000006c6,
      O => blk00000003_sig000006c2
    );
  blk00000003_blk00000576 : MUXCY
    port map (
      CI => blk00000003_sig000006c2,
      DI => blk00000003_sig000006f3,
      S => blk00000003_sig000006c3,
      O => blk00000003_sig000006ef
    );
  blk00000003_blk00000575 : MUXCY
    port map (
      CI => blk00000003_sig000006ef,
      DI => blk00000003_sig000006f1,
      S => blk00000003_sig00000043,
      O => blk00000003_sig000006f2
    );
  blk00000003_blk00000574 : XORCY
    port map (
      CI => blk00000003_sig000006ef,
      LI => blk00000003_sig00000043,
      O => blk00000003_sig000006f0
    );
  blk00000003_blk00000573 : XORCY
    port map (
      CI => blk00000003_sig000006ec,
      LI => blk00000003_sig000006ed,
      O => blk00000003_sig000006ee
    );
  blk00000003_blk00000572 : XORCY
    port map (
      CI => blk00000003_sig000006e9,
      LI => blk00000003_sig000006ea,
      O => blk00000003_sig000006eb
    );
  blk00000003_blk00000571 : XORCY
    port map (
      CI => blk00000003_sig000006e6,
      LI => blk00000003_sig000006e7,
      O => blk00000003_sig000006e8
    );
  blk00000003_blk00000570 : XORCY
    port map (
      CI => blk00000003_sig000006e3,
      LI => blk00000003_sig000006e4,
      O => blk00000003_sig000006e5
    );
  blk00000003_blk0000056f : XORCY
    port map (
      CI => blk00000003_sig000006e0,
      LI => blk00000003_sig000006e1,
      O => blk00000003_sig000006e2
    );
  blk00000003_blk0000056e : XORCY
    port map (
      CI => blk00000003_sig000006dd,
      LI => blk00000003_sig000006de,
      O => blk00000003_sig000006df
    );
  blk00000003_blk0000056d : XORCY
    port map (
      CI => blk00000003_sig000006da,
      LI => blk00000003_sig000006db,
      O => blk00000003_sig000006dc
    );
  blk00000003_blk0000056c : XORCY
    port map (
      CI => blk00000003_sig000006d7,
      LI => blk00000003_sig000006d8,
      O => blk00000003_sig000006d9
    );
  blk00000003_blk0000056b : XORCY
    port map (
      CI => blk00000003_sig000006d4,
      LI => blk00000003_sig000006d5,
      O => blk00000003_sig000006d6
    );
  blk00000003_blk0000056a : XORCY
    port map (
      CI => blk00000003_sig000006d1,
      LI => blk00000003_sig000006d2,
      O => blk00000003_sig000006d3
    );
  blk00000003_blk00000569 : XORCY
    port map (
      CI => blk00000003_sig000006ce,
      LI => blk00000003_sig000006cf,
      O => blk00000003_sig000006d0
    );
  blk00000003_blk00000568 : XORCY
    port map (
      CI => blk00000003_sig000006cb,
      LI => blk00000003_sig000006cc,
      O => blk00000003_sig000006cd
    );
  blk00000003_blk00000567 : XORCY
    port map (
      CI => blk00000003_sig000006c8,
      LI => blk00000003_sig000006c9,
      O => blk00000003_sig000006ca
    );
  blk00000003_blk00000566 : XORCY
    port map (
      CI => blk00000003_sig000006c5,
      LI => blk00000003_sig000006c6,
      O => blk00000003_sig000006c7
    );
  blk00000003_blk00000565 : XORCY
    port map (
      CI => blk00000003_sig000006c2,
      LI => blk00000003_sig000006c3,
      O => blk00000003_sig000006c4
    );
  blk00000003_blk00000564 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000611,
      Q => blk00000003_sig000006c1
    );
  blk00000003_blk00000563 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006b2,
      Q => blk00000003_sig000006c0
    );
  blk00000003_blk00000562 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006b1,
      Q => blk00000003_sig000006bf
    );
  blk00000003_blk00000561 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006b0,
      Q => blk00000003_sig000006be
    );
  blk00000003_blk00000560 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006af,
      Q => blk00000003_sig000006bd
    );
  blk00000003_blk0000055f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ae,
      Q => blk00000003_sig000006bc
    );
  blk00000003_blk0000055e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ad,
      Q => blk00000003_sig000006bb
    );
  blk00000003_blk0000055d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ac,
      Q => blk00000003_sig000006ba
    );
  blk00000003_blk0000055c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ab,
      Q => blk00000003_sig000006b9
    );
  blk00000003_blk0000055b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006aa,
      Q => blk00000003_sig000006b8
    );
  blk00000003_blk0000055a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a9,
      Q => blk00000003_sig000006b7
    );
  blk00000003_blk00000559 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a8,
      Q => blk00000003_sig000006b6
    );
  blk00000003_blk00000558 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a7,
      Q => blk00000003_sig000006b5
    );
  blk00000003_blk00000557 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a6,
      Q => blk00000003_sig000006b4
    );
  blk00000003_blk00000556 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a5,
      Q => blk00000003_sig000006b3
    );
  blk00000003_blk00000555 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000612,
      Q => blk00000003_sig000006b2
    );
  blk00000003_blk00000554 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a4,
      Q => blk00000003_sig000006b1
    );
  blk00000003_blk00000553 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a3,
      Q => blk00000003_sig000006b0
    );
  blk00000003_blk00000552 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a2,
      Q => blk00000003_sig000006af
    );
  blk00000003_blk00000551 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a1,
      Q => blk00000003_sig000006ae
    );
  blk00000003_blk00000550 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a0,
      Q => blk00000003_sig000006ad
    );
  blk00000003_blk0000054f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000069f,
      Q => blk00000003_sig000006ac
    );
  blk00000003_blk0000054e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000069e,
      Q => blk00000003_sig000006ab
    );
  blk00000003_blk0000054d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000069d,
      Q => blk00000003_sig000006aa
    );
  blk00000003_blk0000054c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000069c,
      Q => blk00000003_sig000006a9
    );
  blk00000003_blk0000054b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000069b,
      Q => blk00000003_sig000006a8
    );
  blk00000003_blk0000054a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000069a,
      Q => blk00000003_sig000006a7
    );
  blk00000003_blk00000549 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000699,
      Q => blk00000003_sig000006a6
    );
  blk00000003_blk00000548 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000698,
      Q => blk00000003_sig000006a5
    );
  blk00000003_blk00000547 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000613,
      Q => blk00000003_sig000006a4
    );
  blk00000003_blk00000546 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000697,
      Q => blk00000003_sig000006a3
    );
  blk00000003_blk00000545 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000696,
      Q => blk00000003_sig000006a2
    );
  blk00000003_blk00000544 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000695,
      Q => blk00000003_sig000006a1
    );
  blk00000003_blk00000543 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000694,
      Q => blk00000003_sig000006a0
    );
  blk00000003_blk00000542 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000693,
      Q => blk00000003_sig0000069f
    );
  blk00000003_blk00000541 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000692,
      Q => blk00000003_sig0000069e
    );
  blk00000003_blk00000540 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000691,
      Q => blk00000003_sig0000069d
    );
  blk00000003_blk0000053f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000690,
      Q => blk00000003_sig0000069c
    );
  blk00000003_blk0000053e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000068f,
      Q => blk00000003_sig0000069b
    );
  blk00000003_blk0000053d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000068e,
      Q => blk00000003_sig0000069a
    );
  blk00000003_blk0000053c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000068d,
      Q => blk00000003_sig00000699
    );
  blk00000003_blk0000053b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000068c,
      Q => blk00000003_sig00000698
    );
  blk00000003_blk0000053a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000614,
      Q => blk00000003_sig00000697
    );
  blk00000003_blk00000539 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000068b,
      Q => blk00000003_sig00000696
    );
  blk00000003_blk00000538 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000068a,
      Q => blk00000003_sig00000695
    );
  blk00000003_blk00000537 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000689,
      Q => blk00000003_sig00000694
    );
  blk00000003_blk00000536 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000688,
      Q => blk00000003_sig00000693
    );
  blk00000003_blk00000535 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000687,
      Q => blk00000003_sig00000692
    );
  blk00000003_blk00000534 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000686,
      Q => blk00000003_sig00000691
    );
  blk00000003_blk00000533 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000685,
      Q => blk00000003_sig00000690
    );
  blk00000003_blk00000532 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000684,
      Q => blk00000003_sig0000068f
    );
  blk00000003_blk00000531 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000683,
      Q => blk00000003_sig0000068e
    );
  blk00000003_blk00000530 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000682,
      Q => blk00000003_sig0000068d
    );
  blk00000003_blk0000052f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000681,
      Q => blk00000003_sig0000068c
    );
  blk00000003_blk0000052e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000615,
      Q => blk00000003_sig0000068b
    );
  blk00000003_blk0000052d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000680,
      Q => blk00000003_sig0000068a
    );
  blk00000003_blk0000052c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000067f,
      Q => blk00000003_sig00000689
    );
  blk00000003_blk0000052b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000067e,
      Q => blk00000003_sig00000688
    );
  blk00000003_blk0000052a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000067d,
      Q => blk00000003_sig00000687
    );
  blk00000003_blk00000529 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000067c,
      Q => blk00000003_sig00000686
    );
  blk00000003_blk00000528 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000067b,
      Q => blk00000003_sig00000685
    );
  blk00000003_blk00000527 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000067a,
      Q => blk00000003_sig00000684
    );
  blk00000003_blk00000526 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000679,
      Q => blk00000003_sig00000683
    );
  blk00000003_blk00000525 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000678,
      Q => blk00000003_sig00000682
    );
  blk00000003_blk00000524 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000677,
      Q => blk00000003_sig00000681
    );
  blk00000003_blk00000523 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000616,
      Q => blk00000003_sig00000680
    );
  blk00000003_blk00000522 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000676,
      Q => blk00000003_sig0000067f
    );
  blk00000003_blk00000521 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000675,
      Q => blk00000003_sig0000067e
    );
  blk00000003_blk00000520 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000674,
      Q => blk00000003_sig0000067d
    );
  blk00000003_blk0000051f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000673,
      Q => blk00000003_sig0000067c
    );
  blk00000003_blk0000051e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000672,
      Q => blk00000003_sig0000067b
    );
  blk00000003_blk0000051d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000671,
      Q => blk00000003_sig0000067a
    );
  blk00000003_blk0000051c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000670,
      Q => blk00000003_sig00000679
    );
  blk00000003_blk0000051b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000066f,
      Q => blk00000003_sig00000678
    );
  blk00000003_blk0000051a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000066e,
      Q => blk00000003_sig00000677
    );
  blk00000003_blk00000519 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000617,
      Q => blk00000003_sig00000676
    );
  blk00000003_blk00000518 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000066d,
      Q => blk00000003_sig00000675
    );
  blk00000003_blk00000517 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000066c,
      Q => blk00000003_sig00000674
    );
  blk00000003_blk00000516 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000066b,
      Q => blk00000003_sig00000673
    );
  blk00000003_blk00000515 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000066a,
      Q => blk00000003_sig00000672
    );
  blk00000003_blk00000514 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000669,
      Q => blk00000003_sig00000671
    );
  blk00000003_blk00000513 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000668,
      Q => blk00000003_sig00000670
    );
  blk00000003_blk00000512 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000667,
      Q => blk00000003_sig0000066f
    );
  blk00000003_blk00000511 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000666,
      Q => blk00000003_sig0000066e
    );
  blk00000003_blk00000510 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000618,
      Q => blk00000003_sig0000066d
    );
  blk00000003_blk0000050f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000068,
      Q => blk00000003_sig0000066c
    );
  blk00000003_blk0000050e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006a,
      Q => blk00000003_sig0000066b
    );
  blk00000003_blk0000050d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006c,
      Q => blk00000003_sig0000066a
    );
  blk00000003_blk0000050c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006e,
      Q => blk00000003_sig00000669
    );
  blk00000003_blk0000050b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000070,
      Q => blk00000003_sig00000668
    );
  blk00000003_blk0000050a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000072,
      Q => blk00000003_sig00000667
    );
  blk00000003_blk00000509 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000074,
      Q => blk00000003_sig00000666
    );
  blk00000003_blk00000508 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000665,
      Q => blk00000003_sig0000005f
    );
  blk00000003_blk00000507 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000664,
      Q => blk00000003_sig00000060
    );
  blk00000003_blk00000506 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000663,
      Q => blk00000003_sig00000061
    );
  blk00000003_blk00000505 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000662,
      Q => blk00000003_sig00000062
    );
  blk00000003_blk00000504 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000661,
      Q => blk00000003_sig00000063
    );
  blk00000003_blk00000503 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000660,
      Q => blk00000003_sig00000064
    );
  blk00000003_blk00000502 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000065f,
      Q => blk00000003_sig00000065
    );
  blk00000003_blk00000501 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000065e,
      Q => blk00000003_sig0000041b
    );
  blk00000003_blk00000500 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000065d,
      Q => blk00000003_sig00000665
    );
  blk00000003_blk000004ff : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000065c,
      Q => blk00000003_sig00000664
    );
  blk00000003_blk000004fe : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000065b,
      Q => blk00000003_sig00000663
    );
  blk00000003_blk000004fd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000065a,
      Q => blk00000003_sig00000662
    );
  blk00000003_blk000004fc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000659,
      Q => blk00000003_sig00000661
    );
  blk00000003_blk000004fb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000658,
      Q => blk00000003_sig00000660
    );
  blk00000003_blk000004fa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000657,
      Q => blk00000003_sig0000065f
    );
  blk00000003_blk000004f9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000656,
      Q => blk00000003_sig0000065e
    );
  blk00000003_blk000004f8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000655,
      Q => blk00000003_sig000003d5
    );
  blk00000003_blk000004f7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000654,
      Q => blk00000003_sig0000065d
    );
  blk00000003_blk000004f6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000653,
      Q => blk00000003_sig0000065c
    );
  blk00000003_blk000004f5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000652,
      Q => blk00000003_sig0000065b
    );
  blk00000003_blk000004f4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000651,
      Q => blk00000003_sig0000065a
    );
  blk00000003_blk000004f3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000650,
      Q => blk00000003_sig00000659
    );
  blk00000003_blk000004f2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000064f,
      Q => blk00000003_sig00000658
    );
  blk00000003_blk000004f1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000064e,
      Q => blk00000003_sig00000657
    );
  blk00000003_blk000004f0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000064d,
      Q => blk00000003_sig00000656
    );
  blk00000003_blk000004ef : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000064c,
      Q => blk00000003_sig00000655
    );
  blk00000003_blk000004ee : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000064b,
      Q => blk00000003_sig0000038f
    );
  blk00000003_blk000004ed : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000064a,
      Q => blk00000003_sig00000654
    );
  blk00000003_blk000004ec : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000649,
      Q => blk00000003_sig00000653
    );
  blk00000003_blk000004eb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000648,
      Q => blk00000003_sig00000652
    );
  blk00000003_blk000004ea : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000647,
      Q => blk00000003_sig00000651
    );
  blk00000003_blk000004e9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000646,
      Q => blk00000003_sig00000650
    );
  blk00000003_blk000004e8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000645,
      Q => blk00000003_sig0000064f
    );
  blk00000003_blk000004e7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000644,
      Q => blk00000003_sig0000064e
    );
  blk00000003_blk000004e6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000643,
      Q => blk00000003_sig0000064d
    );
  blk00000003_blk000004e5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000642,
      Q => blk00000003_sig0000064c
    );
  blk00000003_blk000004e4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000641,
      Q => blk00000003_sig0000064b
    );
  blk00000003_blk000004e3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000640,
      Q => blk00000003_sig00000349
    );
  blk00000003_blk000004e2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000063f,
      Q => blk00000003_sig0000064a
    );
  blk00000003_blk000004e1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000063e,
      Q => blk00000003_sig00000649
    );
  blk00000003_blk000004e0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000063d,
      Q => blk00000003_sig00000648
    );
  blk00000003_blk000004df : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000063c,
      Q => blk00000003_sig00000647
    );
  blk00000003_blk000004de : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000063b,
      Q => blk00000003_sig00000646
    );
  blk00000003_blk000004dd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000063a,
      Q => blk00000003_sig00000645
    );
  blk00000003_blk000004dc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000639,
      Q => blk00000003_sig00000644
    );
  blk00000003_blk000004db : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000638,
      Q => blk00000003_sig00000643
    );
  blk00000003_blk000004da : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000637,
      Q => blk00000003_sig00000642
    );
  blk00000003_blk000004d9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000636,
      Q => blk00000003_sig00000641
    );
  blk00000003_blk000004d8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000635,
      Q => blk00000003_sig00000640
    );
  blk00000003_blk000004d7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000634,
      Q => blk00000003_sig00000303
    );
  blk00000003_blk000004d6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000633,
      Q => blk00000003_sig0000063f
    );
  blk00000003_blk000004d5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000632,
      Q => blk00000003_sig0000063e
    );
  blk00000003_blk000004d4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000631,
      Q => blk00000003_sig0000063d
    );
  blk00000003_blk000004d3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000630,
      Q => blk00000003_sig0000063c
    );
  blk00000003_blk000004d2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000062f,
      Q => blk00000003_sig0000063b
    );
  blk00000003_blk000004d1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000062e,
      Q => blk00000003_sig0000063a
    );
  blk00000003_blk000004d0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000062d,
      Q => blk00000003_sig00000639
    );
  blk00000003_blk000004cf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000062c,
      Q => blk00000003_sig00000638
    );
  blk00000003_blk000004ce : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000062b,
      Q => blk00000003_sig00000637
    );
  blk00000003_blk000004cd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000062a,
      Q => blk00000003_sig00000636
    );
  blk00000003_blk000004cc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000629,
      Q => blk00000003_sig00000635
    );
  blk00000003_blk000004cb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000628,
      Q => blk00000003_sig00000634
    );
  blk00000003_blk000004ca : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000627,
      Q => blk00000003_sig000002bd
    );
  blk00000003_blk000004c9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000626,
      Q => blk00000003_sig00000633
    );
  blk00000003_blk000004c8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000625,
      Q => blk00000003_sig00000632
    );
  blk00000003_blk000004c7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000624,
      Q => blk00000003_sig00000631
    );
  blk00000003_blk000004c6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000623,
      Q => blk00000003_sig00000630
    );
  blk00000003_blk000004c5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000622,
      Q => blk00000003_sig0000062f
    );
  blk00000003_blk000004c4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000621,
      Q => blk00000003_sig0000062e
    );
  blk00000003_blk000004c3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000620,
      Q => blk00000003_sig0000062d
    );
  blk00000003_blk000004c2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000061f,
      Q => blk00000003_sig0000062c
    );
  blk00000003_blk000004c1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000061e,
      Q => blk00000003_sig0000062b
    );
  blk00000003_blk000004c0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000061d,
      Q => blk00000003_sig0000062a
    );
  blk00000003_blk000004bf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000061c,
      Q => blk00000003_sig00000629
    );
  blk00000003_blk000004be : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000061b,
      Q => blk00000003_sig00000628
    );
  blk00000003_blk000004bd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000061a,
      Q => blk00000003_sig00000627
    );
  blk00000003_blk000004bc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000619,
      Q => blk00000003_sig00000277
    );
  blk00000003_blk000004bb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000aa,
      Q => blk00000003_sig00000626
    );
  blk00000003_blk000004ba : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a9,
      Q => blk00000003_sig00000625
    );
  blk00000003_blk000004b9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a8,
      Q => blk00000003_sig00000624
    );
  blk00000003_blk000004b8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a7,
      Q => blk00000003_sig00000623
    );
  blk00000003_blk000004b7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a6,
      Q => blk00000003_sig00000622
    );
  blk00000003_blk000004b6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a5,
      Q => blk00000003_sig00000621
    );
  blk00000003_blk000004b5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a4,
      Q => blk00000003_sig00000620
    );
  blk00000003_blk000004b4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a3,
      Q => blk00000003_sig0000061f
    );
  blk00000003_blk000004b3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a2,
      Q => blk00000003_sig0000061e
    );
  blk00000003_blk000004b2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a1,
      Q => blk00000003_sig0000061d
    );
  blk00000003_blk000004b1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a0,
      Q => blk00000003_sig0000061c
    );
  blk00000003_blk000004b0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000009f,
      Q => blk00000003_sig0000061b
    );
  blk00000003_blk000004af : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000009e,
      Q => blk00000003_sig0000061a
    );
  blk00000003_blk000004ae : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000009d,
      Q => blk00000003_sig00000619
    );
  blk00000003_blk000004ad : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000009c,
      Q => blk00000003_sig00000231
    );
  blk00000003_blk000004ac : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001eb,
      Q => blk00000003_sig0000022b
    );
  blk00000003_blk000004ab : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001e8,
      Q => blk00000003_sig0000022a
    );
  blk00000003_blk000004aa : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001e5,
      Q => blk00000003_sig00000229
    );
  blk00000003_blk000004a9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001e2,
      Q => blk00000003_sig00000228
    );
  blk00000003_blk000004a8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001df,
      Q => blk00000003_sig00000227
    );
  blk00000003_blk000004a7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001dc,
      Q => blk00000003_sig00000226
    );
  blk00000003_blk000004a6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001d9,
      Q => blk00000003_sig00000225
    );
  blk00000003_blk000004a5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001d6,
      Q => blk00000003_sig00000224
    );
  blk00000003_blk000004a4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001d3,
      Q => blk00000003_sig00000223
    );
  blk00000003_blk000004a3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001d0,
      Q => blk00000003_sig00000222
    );
  blk00000003_blk000004a2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001cd,
      Q => blk00000003_sig00000221
    );
  blk00000003_blk000004a1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001ca,
      Q => blk00000003_sig00000220
    );
  blk00000003_blk000004a0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001c7,
      Q => blk00000003_sig0000021f
    );
  blk00000003_blk0000049f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001c4,
      Q => blk00000003_sig0000021e
    );
  blk00000003_blk0000049e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001c1,
      Q => blk00000003_sig0000021d
    );
  blk00000003_blk0000049d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001be,
      Q => blk00000003_sig0000022c
    );
  blk00000003_blk0000049c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000230,
      Q => blk00000003_sig00000271
    );
  blk00000003_blk0000049b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000021c,
      Q => blk00000003_sig00000270
    );
  blk00000003_blk0000049a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000219,
      Q => blk00000003_sig0000026f
    );
  blk00000003_blk00000499 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000216,
      Q => blk00000003_sig0000026e
    );
  blk00000003_blk00000498 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000213,
      Q => blk00000003_sig0000026d
    );
  blk00000003_blk00000497 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000210,
      Q => blk00000003_sig0000026c
    );
  blk00000003_blk00000496 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000020d,
      Q => blk00000003_sig0000026b
    );
  blk00000003_blk00000495 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000020a,
      Q => blk00000003_sig0000026a
    );
  blk00000003_blk00000494 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000207,
      Q => blk00000003_sig00000269
    );
  blk00000003_blk00000493 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000204,
      Q => blk00000003_sig00000268
    );
  blk00000003_blk00000492 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000201,
      Q => blk00000003_sig00000267
    );
  blk00000003_blk00000491 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001fe,
      Q => blk00000003_sig00000266
    );
  blk00000003_blk00000490 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001fb,
      Q => blk00000003_sig00000265
    );
  blk00000003_blk0000048f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001f8,
      Q => blk00000003_sig00000264
    );
  blk00000003_blk0000048e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001f5,
      Q => blk00000003_sig00000263
    );
  blk00000003_blk0000048d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001f2,
      Q => blk00000003_sig00000272
    );
  blk00000003_blk0000048c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001ef,
      Q => blk00000003_sig00000087
    );
  blk00000003_blk0000048b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000276,
      Q => blk00000003_sig000002b7
    );
  blk00000003_blk0000048a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000262,
      Q => blk00000003_sig000002b6
    );
  blk00000003_blk00000489 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000025f,
      Q => blk00000003_sig000002b5
    );
  blk00000003_blk00000488 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000025c,
      Q => blk00000003_sig000002b4
    );
  blk00000003_blk00000487 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000259,
      Q => blk00000003_sig000002b3
    );
  blk00000003_blk00000486 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000256,
      Q => blk00000003_sig000002b2
    );
  blk00000003_blk00000485 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000253,
      Q => blk00000003_sig000002b1
    );
  blk00000003_blk00000484 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000250,
      Q => blk00000003_sig000002b0
    );
  blk00000003_blk00000483 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000024d,
      Q => blk00000003_sig000002af
    );
  blk00000003_blk00000482 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000024a,
      Q => blk00000003_sig000002ae
    );
  blk00000003_blk00000481 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000247,
      Q => blk00000003_sig000002ad
    );
  blk00000003_blk00000480 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000244,
      Q => blk00000003_sig000002ac
    );
  blk00000003_blk0000047f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000241,
      Q => blk00000003_sig000002ab
    );
  blk00000003_blk0000047e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000023e,
      Q => blk00000003_sig000002aa
    );
  blk00000003_blk0000047d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000023b,
      Q => blk00000003_sig000002a9
    );
  blk00000003_blk0000047c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000238,
      Q => blk00000003_sig000002b8
    );
  blk00000003_blk0000047b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000235,
      Q => blk00000003_sig00000084
    );
  blk00000003_blk0000047a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002bc,
      Q => blk00000003_sig000002fd
    );
  blk00000003_blk00000479 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002a8,
      Q => blk00000003_sig000002fc
    );
  blk00000003_blk00000478 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002a5,
      Q => blk00000003_sig000002fb
    );
  blk00000003_blk00000477 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002a2,
      Q => blk00000003_sig000002fa
    );
  blk00000003_blk00000476 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000029f,
      Q => blk00000003_sig000002f9
    );
  blk00000003_blk00000475 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000029c,
      Q => blk00000003_sig000002f8
    );
  blk00000003_blk00000474 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000299,
      Q => blk00000003_sig000002f7
    );
  blk00000003_blk00000473 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000296,
      Q => blk00000003_sig000002f6
    );
  blk00000003_blk00000472 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000293,
      Q => blk00000003_sig000002f5
    );
  blk00000003_blk00000471 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000290,
      Q => blk00000003_sig000002f4
    );
  blk00000003_blk00000470 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000028d,
      Q => blk00000003_sig000002f3
    );
  blk00000003_blk0000046f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000028a,
      Q => blk00000003_sig000002f2
    );
  blk00000003_blk0000046e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000287,
      Q => blk00000003_sig000002f1
    );
  blk00000003_blk0000046d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000284,
      Q => blk00000003_sig000002f0
    );
  blk00000003_blk0000046c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000281,
      Q => blk00000003_sig000002ef
    );
  blk00000003_blk0000046b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000027e,
      Q => blk00000003_sig000002fe
    );
  blk00000003_blk0000046a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000027b,
      Q => blk00000003_sig00000080
    );
  blk00000003_blk00000469 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000302,
      Q => blk00000003_sig00000343
    );
  blk00000003_blk00000468 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002ee,
      Q => blk00000003_sig00000342
    );
  blk00000003_blk00000467 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002eb,
      Q => blk00000003_sig00000341
    );
  blk00000003_blk00000466 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002e8,
      Q => blk00000003_sig00000340
    );
  blk00000003_blk00000465 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002e5,
      Q => blk00000003_sig0000033f
    );
  blk00000003_blk00000464 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002e2,
      Q => blk00000003_sig0000033e
    );
  blk00000003_blk00000463 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002df,
      Q => blk00000003_sig0000033d
    );
  blk00000003_blk00000462 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002dc,
      Q => blk00000003_sig0000033c
    );
  blk00000003_blk00000461 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002d9,
      Q => blk00000003_sig0000033b
    );
  blk00000003_blk00000460 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002d6,
      Q => blk00000003_sig0000033a
    );
  blk00000003_blk0000045f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002d3,
      Q => blk00000003_sig00000339
    );
  blk00000003_blk0000045e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002d0,
      Q => blk00000003_sig00000338
    );
  blk00000003_blk0000045d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002cd,
      Q => blk00000003_sig00000337
    );
  blk00000003_blk0000045c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002ca,
      Q => blk00000003_sig00000336
    );
  blk00000003_blk0000045b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002c7,
      Q => blk00000003_sig00000335
    );
  blk00000003_blk0000045a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002c4,
      Q => blk00000003_sig00000344
    );
  blk00000003_blk00000459 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002c1,
      Q => blk00000003_sig0000007b
    );
  blk00000003_blk00000458 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000348,
      Q => blk00000003_sig00000389
    );
  blk00000003_blk00000457 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000334,
      Q => blk00000003_sig00000388
    );
  blk00000003_blk00000456 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000331,
      Q => blk00000003_sig00000387
    );
  blk00000003_blk00000455 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000032e,
      Q => blk00000003_sig00000386
    );
  blk00000003_blk00000454 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000032b,
      Q => blk00000003_sig00000385
    );
  blk00000003_blk00000453 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000328,
      Q => blk00000003_sig00000384
    );
  blk00000003_blk00000452 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000325,
      Q => blk00000003_sig00000383
    );
  blk00000003_blk00000451 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000322,
      Q => blk00000003_sig00000382
    );
  blk00000003_blk00000450 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000031f,
      Q => blk00000003_sig00000381
    );
  blk00000003_blk0000044f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000031c,
      Q => blk00000003_sig00000380
    );
  blk00000003_blk0000044e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000319,
      Q => blk00000003_sig0000037f
    );
  blk00000003_blk0000044d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000316,
      Q => blk00000003_sig0000037e
    );
  blk00000003_blk0000044c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000313,
      Q => blk00000003_sig0000037d
    );
  blk00000003_blk0000044b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000310,
      Q => blk00000003_sig0000037c
    );
  blk00000003_blk0000044a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000030d,
      Q => blk00000003_sig0000037b
    );
  blk00000003_blk00000449 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000030a,
      Q => blk00000003_sig0000038a
    );
  blk00000003_blk00000448 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000307,
      Q => blk00000003_sig00000075
    );
  blk00000003_blk00000447 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000038e,
      Q => blk00000003_sig000003cf
    );
  blk00000003_blk00000446 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000037a,
      Q => blk00000003_sig000003ce
    );
  blk00000003_blk00000445 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000377,
      Q => blk00000003_sig000003cd
    );
  blk00000003_blk00000444 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000374,
      Q => blk00000003_sig000003cc
    );
  blk00000003_blk00000443 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000371,
      Q => blk00000003_sig000003cb
    );
  blk00000003_blk00000442 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000036e,
      Q => blk00000003_sig000003ca
    );
  blk00000003_blk00000441 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000036b,
      Q => blk00000003_sig000003c9
    );
  blk00000003_blk00000440 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000368,
      Q => blk00000003_sig000003c8
    );
  blk00000003_blk0000043f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000365,
      Q => blk00000003_sig000003c7
    );
  blk00000003_blk0000043e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000362,
      Q => blk00000003_sig000003c6
    );
  blk00000003_blk0000043d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000035f,
      Q => blk00000003_sig000003c5
    );
  blk00000003_blk0000043c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000035c,
      Q => blk00000003_sig000003c4
    );
  blk00000003_blk0000043b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000359,
      Q => blk00000003_sig000003c3
    );
  blk00000003_blk0000043a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000356,
      Q => blk00000003_sig000003c2
    );
  blk00000003_blk00000439 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000353,
      Q => blk00000003_sig000003c1
    );
  blk00000003_blk00000438 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000350,
      Q => blk00000003_sig000003d0
    );
  blk00000003_blk00000437 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000034d,
      Q => blk00000003_sig00000067
    );
  blk00000003_blk00000436 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003d4,
      Q => blk00000003_sig00000415
    );
  blk00000003_blk00000435 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003c0,
      Q => blk00000003_sig00000414
    );
  blk00000003_blk00000434 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003bd,
      Q => blk00000003_sig00000413
    );
  blk00000003_blk00000433 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003ba,
      Q => blk00000003_sig00000412
    );
  blk00000003_blk00000432 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003b7,
      Q => blk00000003_sig00000411
    );
  blk00000003_blk00000431 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003b4,
      Q => blk00000003_sig00000410
    );
  blk00000003_blk00000430 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003b1,
      Q => blk00000003_sig0000040f
    );
  blk00000003_blk0000042f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003ae,
      Q => blk00000003_sig0000040e
    );
  blk00000003_blk0000042e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003ab,
      Q => blk00000003_sig0000040d
    );
  blk00000003_blk0000042d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003a8,
      Q => blk00000003_sig0000040c
    );
  blk00000003_blk0000042c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003a5,
      Q => blk00000003_sig0000040b
    );
  blk00000003_blk0000042b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003a2,
      Q => blk00000003_sig0000040a
    );
  blk00000003_blk0000042a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000039f,
      Q => blk00000003_sig00000409
    );
  blk00000003_blk00000429 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000039c,
      Q => blk00000003_sig00000408
    );
  blk00000003_blk00000428 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000399,
      Q => blk00000003_sig00000407
    );
  blk00000003_blk00000427 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000396,
      Q => blk00000003_sig00000416
    );
  blk00000003_blk00000426 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000393,
      Q => blk00000003_sig00000618
    );
  blk00000003_blk00000425 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000041a,
      Q => blk00000003_sig0000045b
    );
  blk00000003_blk00000424 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000406,
      Q => blk00000003_sig0000045a
    );
  blk00000003_blk00000423 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000403,
      Q => blk00000003_sig00000459
    );
  blk00000003_blk00000422 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000400,
      Q => blk00000003_sig00000458
    );
  blk00000003_blk00000421 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003fd,
      Q => blk00000003_sig00000457
    );
  blk00000003_blk00000420 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003fa,
      Q => blk00000003_sig00000456
    );
  blk00000003_blk0000041f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003f7,
      Q => blk00000003_sig00000455
    );
  blk00000003_blk0000041e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003f4,
      Q => blk00000003_sig00000454
    );
  blk00000003_blk0000041d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003f1,
      Q => blk00000003_sig00000453
    );
  blk00000003_blk0000041c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003ee,
      Q => blk00000003_sig00000452
    );
  blk00000003_blk0000041b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003eb,
      Q => blk00000003_sig00000451
    );
  blk00000003_blk0000041a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003e8,
      Q => blk00000003_sig00000450
    );
  blk00000003_blk00000419 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003e5,
      Q => blk00000003_sig0000044f
    );
  blk00000003_blk00000418 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003e2,
      Q => blk00000003_sig0000044e
    );
  blk00000003_blk00000417 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003df,
      Q => blk00000003_sig0000044d
    );
  blk00000003_blk00000416 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003dc,
      Q => blk00000003_sig0000045c
    );
  blk00000003_blk00000415 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003d9,
      Q => blk00000003_sig00000617
    );
  blk00000003_blk00000414 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000460,
      Q => blk00000003_sig000004a0
    );
  blk00000003_blk00000413 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000044c,
      Q => blk00000003_sig0000049f
    );
  blk00000003_blk00000412 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000449,
      Q => blk00000003_sig0000049e
    );
  blk00000003_blk00000411 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000446,
      Q => blk00000003_sig0000049d
    );
  blk00000003_blk00000410 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000443,
      Q => blk00000003_sig0000049c
    );
  blk00000003_blk0000040f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000440,
      Q => blk00000003_sig0000049b
    );
  blk00000003_blk0000040e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000043d,
      Q => blk00000003_sig0000049a
    );
  blk00000003_blk0000040d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000043a,
      Q => blk00000003_sig00000499
    );
  blk00000003_blk0000040c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000437,
      Q => blk00000003_sig00000498
    );
  blk00000003_blk0000040b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000434,
      Q => blk00000003_sig00000497
    );
  blk00000003_blk0000040a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000431,
      Q => blk00000003_sig00000496
    );
  blk00000003_blk00000409 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000042e,
      Q => blk00000003_sig00000495
    );
  blk00000003_blk00000408 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000042b,
      Q => blk00000003_sig00000494
    );
  blk00000003_blk00000407 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000428,
      Q => blk00000003_sig00000493
    );
  blk00000003_blk00000406 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000425,
      Q => blk00000003_sig00000492
    );
  blk00000003_blk00000405 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000422,
      Q => blk00000003_sig000004a1
    );
  blk00000003_blk00000404 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000041f,
      Q => blk00000003_sig00000616
    );
  blk00000003_blk00000403 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004a5,
      Q => blk00000003_sig000004e5
    );
  blk00000003_blk00000402 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000491,
      Q => blk00000003_sig000004e4
    );
  blk00000003_blk00000401 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000048e,
      Q => blk00000003_sig000004e3
    );
  blk00000003_blk00000400 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000048b,
      Q => blk00000003_sig000004e2
    );
  blk00000003_blk000003ff : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000488,
      Q => blk00000003_sig000004e1
    );
  blk00000003_blk000003fe : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000485,
      Q => blk00000003_sig000004e0
    );
  blk00000003_blk000003fd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000482,
      Q => blk00000003_sig000004df
    );
  blk00000003_blk000003fc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000047f,
      Q => blk00000003_sig000004de
    );
  blk00000003_blk000003fb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000047c,
      Q => blk00000003_sig000004dd
    );
  blk00000003_blk000003fa : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000479,
      Q => blk00000003_sig000004dc
    );
  blk00000003_blk000003f9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000476,
      Q => blk00000003_sig000004db
    );
  blk00000003_blk000003f8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000473,
      Q => blk00000003_sig000004da
    );
  blk00000003_blk000003f7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000470,
      Q => blk00000003_sig000004d9
    );
  blk00000003_blk000003f6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000046d,
      Q => blk00000003_sig000004d8
    );
  blk00000003_blk000003f5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000046a,
      Q => blk00000003_sig000004d7
    );
  blk00000003_blk000003f4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000467,
      Q => blk00000003_sig000004e6
    );
  blk00000003_blk000003f3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000464,
      Q => blk00000003_sig00000615
    );
  blk00000003_blk000003f2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004ea,
      Q => blk00000003_sig0000052a
    );
  blk00000003_blk000003f1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004d6,
      Q => blk00000003_sig00000529
    );
  blk00000003_blk000003f0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004d3,
      Q => blk00000003_sig00000528
    );
  blk00000003_blk000003ef : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004d0,
      Q => blk00000003_sig00000527
    );
  blk00000003_blk000003ee : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004cd,
      Q => blk00000003_sig00000526
    );
  blk00000003_blk000003ed : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004ca,
      Q => blk00000003_sig00000525
    );
  blk00000003_blk000003ec : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004c7,
      Q => blk00000003_sig00000524
    );
  blk00000003_blk000003eb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004c4,
      Q => blk00000003_sig00000523
    );
  blk00000003_blk000003ea : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004c1,
      Q => blk00000003_sig00000522
    );
  blk00000003_blk000003e9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004be,
      Q => blk00000003_sig00000521
    );
  blk00000003_blk000003e8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004bb,
      Q => blk00000003_sig00000520
    );
  blk00000003_blk000003e7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004b8,
      Q => blk00000003_sig0000051f
    );
  blk00000003_blk000003e6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004b5,
      Q => blk00000003_sig0000051e
    );
  blk00000003_blk000003e5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004b2,
      Q => blk00000003_sig0000051d
    );
  blk00000003_blk000003e4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004af,
      Q => blk00000003_sig0000051c
    );
  blk00000003_blk000003e3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004ac,
      Q => blk00000003_sig0000052b
    );
  blk00000003_blk000003e2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004a9,
      Q => blk00000003_sig00000614
    );
  blk00000003_blk000003e1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000052f,
      Q => blk00000003_sig0000056f
    );
  blk00000003_blk000003e0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000051b,
      Q => blk00000003_sig0000056e
    );
  blk00000003_blk000003df : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000518,
      Q => blk00000003_sig0000056d
    );
  blk00000003_blk000003de : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000515,
      Q => blk00000003_sig0000056c
    );
  blk00000003_blk000003dd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000512,
      Q => blk00000003_sig0000056b
    );
  blk00000003_blk000003dc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000050f,
      Q => blk00000003_sig0000056a
    );
  blk00000003_blk000003db : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000050c,
      Q => blk00000003_sig00000569
    );
  blk00000003_blk000003da : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000509,
      Q => blk00000003_sig00000568
    );
  blk00000003_blk000003d9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000506,
      Q => blk00000003_sig00000567
    );
  blk00000003_blk000003d8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000503,
      Q => blk00000003_sig00000566
    );
  blk00000003_blk000003d7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000500,
      Q => blk00000003_sig00000565
    );
  blk00000003_blk000003d6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004fd,
      Q => blk00000003_sig00000564
    );
  blk00000003_blk000003d5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004fa,
      Q => blk00000003_sig00000563
    );
  blk00000003_blk000003d4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004f7,
      Q => blk00000003_sig00000562
    );
  blk00000003_blk000003d3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004f4,
      Q => blk00000003_sig00000561
    );
  blk00000003_blk000003d2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004f1,
      Q => blk00000003_sig00000570
    );
  blk00000003_blk000003d1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004ee,
      Q => blk00000003_sig00000613
    );
  blk00000003_blk000003d0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000574,
      Q => blk00000003_sig000005b4
    );
  blk00000003_blk000003cf : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000560,
      Q => blk00000003_sig000005b3
    );
  blk00000003_blk000003ce : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000055d,
      Q => blk00000003_sig000005b2
    );
  blk00000003_blk000003cd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000055a,
      Q => blk00000003_sig000005b1
    );
  blk00000003_blk000003cc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000557,
      Q => blk00000003_sig000005b0
    );
  blk00000003_blk000003cb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000554,
      Q => blk00000003_sig000005af
    );
  blk00000003_blk000003ca : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000551,
      Q => blk00000003_sig000005ae
    );
  blk00000003_blk000003c9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000054e,
      Q => blk00000003_sig000005ad
    );
  blk00000003_blk000003c8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000054b,
      Q => blk00000003_sig000005ac
    );
  blk00000003_blk000003c7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000548,
      Q => blk00000003_sig000005ab
    );
  blk00000003_blk000003c6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000545,
      Q => blk00000003_sig000005aa
    );
  blk00000003_blk000003c5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000542,
      Q => blk00000003_sig000005a9
    );
  blk00000003_blk000003c4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000053f,
      Q => blk00000003_sig000005a8
    );
  blk00000003_blk000003c3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000053c,
      Q => blk00000003_sig000005a7
    );
  blk00000003_blk000003c2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000539,
      Q => blk00000003_sig000005a6
    );
  blk00000003_blk000003c1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000536,
      Q => blk00000003_sig000005b5
    );
  blk00000003_blk000003c0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000533,
      Q => blk00000003_sig00000612
    );
  blk00000003_blk000003bf : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005b9,
      Q => blk00000003_sig000005f9
    );
  blk00000003_blk000003be : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005a5,
      Q => blk00000003_sig000005f8
    );
  blk00000003_blk000003bd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005a2,
      Q => blk00000003_sig000005f7
    );
  blk00000003_blk000003bc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000059f,
      Q => blk00000003_sig000005f6
    );
  blk00000003_blk000003bb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000059c,
      Q => blk00000003_sig000005f5
    );
  blk00000003_blk000003ba : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000599,
      Q => blk00000003_sig000005f4
    );
  blk00000003_blk000003b9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000596,
      Q => blk00000003_sig000005f3
    );
  blk00000003_blk000003b8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000593,
      Q => blk00000003_sig000005f2
    );
  blk00000003_blk000003b7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000590,
      Q => blk00000003_sig000005f1
    );
  blk00000003_blk000003b6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000058d,
      Q => blk00000003_sig000005f0
    );
  blk00000003_blk000003b5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000058a,
      Q => blk00000003_sig000005ef
    );
  blk00000003_blk000003b4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000587,
      Q => blk00000003_sig000005ee
    );
  blk00000003_blk000003b3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000584,
      Q => blk00000003_sig000005ed
    );
  blk00000003_blk000003b2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000581,
      Q => blk00000003_sig000005ec
    );
  blk00000003_blk000003b1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000057e,
      Q => blk00000003_sig000005eb
    );
  blk00000003_blk000003b0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000057b,
      Q => blk00000003_sig000005fa
    );
  blk00000003_blk000003af : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000578,
      Q => blk00000003_sig00000611
    );
  blk00000003_blk000003ae : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005fe,
      Q => blk00000003_sig00000610
    );
  blk00000003_blk000003ad : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005ea,
      Q => blk00000003_sig0000060f
    );
  blk00000003_blk000003ac : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005e7,
      Q => blk00000003_sig0000060e
    );
  blk00000003_blk000003ab : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005e4,
      Q => blk00000003_sig0000060d
    );
  blk00000003_blk000003aa : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005e1,
      Q => blk00000003_sig0000060c
    );
  blk00000003_blk000003a9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005de,
      Q => blk00000003_sig0000060b
    );
  blk00000003_blk000003a8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005db,
      Q => blk00000003_sig0000060a
    );
  blk00000003_blk000003a7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005d8,
      Q => blk00000003_sig00000609
    );
  blk00000003_blk000003a6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005d5,
      Q => blk00000003_sig00000608
    );
  blk00000003_blk000003a5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005d2,
      Q => blk00000003_sig00000607
    );
  blk00000003_blk000003a4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005cf,
      Q => blk00000003_sig00000606
    );
  blk00000003_blk000003a3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005cc,
      Q => blk00000003_sig00000605
    );
  blk00000003_blk000003a2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005c9,
      Q => blk00000003_sig00000604
    );
  blk00000003_blk000003a1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005c6,
      Q => blk00000003_sig00000603
    );
  blk00000003_blk000003a0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005c3,
      Q => blk00000003_sig00000602
    );
  blk00000003_blk0000039f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005c0,
      Q => blk00000003_sig00000601
    );
  blk00000003_blk0000039e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005bd,
      Q => blk00000003_sig00000600
    );
  blk00000003_blk0000039d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005fb,
      Q => blk00000003_sig000005ff
    );
  blk00000003_blk0000039c : MUXCY
    port map (
      CI => blk00000003_sig000005fc,
      DI => blk00000003_sig0000008a,
      S => blk00000003_sig000005fd,
      O => blk00000003_sig000005e8
    );
  blk00000003_blk0000039b : XORCY
    port map (
      CI => blk00000003_sig000005fc,
      LI => blk00000003_sig000005fd,
      O => blk00000003_sig000005fe
    );
  blk00000003_blk0000039a : MUXCY
    port map (
      CI => blk00000003_sig000005bb,
      DI => blk00000003_sig000005fa,
      S => blk00000003_sig000005bc,
      O => blk00000003_sig000005fb
    );
  blk00000003_blk00000399 : MUXCY
    port map (
      CI => blk00000003_sig000005e8,
      DI => blk00000003_sig000005f9,
      S => blk00000003_sig000005e9,
      O => blk00000003_sig000005e5
    );
  blk00000003_blk00000398 : MUXCY
    port map (
      CI => blk00000003_sig000005e5,
      DI => blk00000003_sig000005f8,
      S => blk00000003_sig000005e6,
      O => blk00000003_sig000005e2
    );
  blk00000003_blk00000397 : MUXCY
    port map (
      CI => blk00000003_sig000005e2,
      DI => blk00000003_sig000005f7,
      S => blk00000003_sig000005e3,
      O => blk00000003_sig000005df
    );
  blk00000003_blk00000396 : MUXCY
    port map (
      CI => blk00000003_sig000005df,
      DI => blk00000003_sig000005f6,
      S => blk00000003_sig000005e0,
      O => blk00000003_sig000005dc
    );
  blk00000003_blk00000395 : MUXCY
    port map (
      CI => blk00000003_sig000005dc,
      DI => blk00000003_sig000005f5,
      S => blk00000003_sig000005dd,
      O => blk00000003_sig000005d9
    );
  blk00000003_blk00000394 : MUXCY
    port map (
      CI => blk00000003_sig000005d9,
      DI => blk00000003_sig000005f4,
      S => blk00000003_sig000005da,
      O => blk00000003_sig000005d6
    );
  blk00000003_blk00000393 : MUXCY
    port map (
      CI => blk00000003_sig000005d6,
      DI => blk00000003_sig000005f3,
      S => blk00000003_sig000005d7,
      O => blk00000003_sig000005d3
    );
  blk00000003_blk00000392 : MUXCY
    port map (
      CI => blk00000003_sig000005d3,
      DI => blk00000003_sig000005f2,
      S => blk00000003_sig000005d4,
      O => blk00000003_sig000005d0
    );
  blk00000003_blk00000391 : MUXCY
    port map (
      CI => blk00000003_sig000005d0,
      DI => blk00000003_sig000005f1,
      S => blk00000003_sig000005d1,
      O => blk00000003_sig000005cd
    );
  blk00000003_blk00000390 : MUXCY
    port map (
      CI => blk00000003_sig000005cd,
      DI => blk00000003_sig000005f0,
      S => blk00000003_sig000005ce,
      O => blk00000003_sig000005ca
    );
  blk00000003_blk0000038f : MUXCY
    port map (
      CI => blk00000003_sig000005ca,
      DI => blk00000003_sig000005ef,
      S => blk00000003_sig000005cb,
      O => blk00000003_sig000005c7
    );
  blk00000003_blk0000038e : MUXCY
    port map (
      CI => blk00000003_sig000005c7,
      DI => blk00000003_sig000005ee,
      S => blk00000003_sig000005c8,
      O => blk00000003_sig000005c4
    );
  blk00000003_blk0000038d : MUXCY
    port map (
      CI => blk00000003_sig000005c4,
      DI => blk00000003_sig000005ed,
      S => blk00000003_sig000005c5,
      O => blk00000003_sig000005c1
    );
  blk00000003_blk0000038c : MUXCY
    port map (
      CI => blk00000003_sig000005c1,
      DI => blk00000003_sig000005ec,
      S => blk00000003_sig000005c2,
      O => blk00000003_sig000005be
    );
  blk00000003_blk0000038b : MUXCY
    port map (
      CI => blk00000003_sig000005be,
      DI => blk00000003_sig000005eb,
      S => blk00000003_sig000005bf,
      O => blk00000003_sig000005bb
    );
  blk00000003_blk0000038a : XORCY
    port map (
      CI => blk00000003_sig000005e8,
      LI => blk00000003_sig000005e9,
      O => blk00000003_sig000005ea
    );
  blk00000003_blk00000389 : XORCY
    port map (
      CI => blk00000003_sig000005e5,
      LI => blk00000003_sig000005e6,
      O => blk00000003_sig000005e7
    );
  blk00000003_blk00000388 : XORCY
    port map (
      CI => blk00000003_sig000005e2,
      LI => blk00000003_sig000005e3,
      O => blk00000003_sig000005e4
    );
  blk00000003_blk00000387 : XORCY
    port map (
      CI => blk00000003_sig000005df,
      LI => blk00000003_sig000005e0,
      O => blk00000003_sig000005e1
    );
  blk00000003_blk00000386 : XORCY
    port map (
      CI => blk00000003_sig000005dc,
      LI => blk00000003_sig000005dd,
      O => blk00000003_sig000005de
    );
  blk00000003_blk00000385 : XORCY
    port map (
      CI => blk00000003_sig000005d9,
      LI => blk00000003_sig000005da,
      O => blk00000003_sig000005db
    );
  blk00000003_blk00000384 : XORCY
    port map (
      CI => blk00000003_sig000005d6,
      LI => blk00000003_sig000005d7,
      O => blk00000003_sig000005d8
    );
  blk00000003_blk00000383 : XORCY
    port map (
      CI => blk00000003_sig000005d3,
      LI => blk00000003_sig000005d4,
      O => blk00000003_sig000005d5
    );
  blk00000003_blk00000382 : XORCY
    port map (
      CI => blk00000003_sig000005d0,
      LI => blk00000003_sig000005d1,
      O => blk00000003_sig000005d2
    );
  blk00000003_blk00000381 : XORCY
    port map (
      CI => blk00000003_sig000005cd,
      LI => blk00000003_sig000005ce,
      O => blk00000003_sig000005cf
    );
  blk00000003_blk00000380 : XORCY
    port map (
      CI => blk00000003_sig000005ca,
      LI => blk00000003_sig000005cb,
      O => blk00000003_sig000005cc
    );
  blk00000003_blk0000037f : XORCY
    port map (
      CI => blk00000003_sig000005c7,
      LI => blk00000003_sig000005c8,
      O => blk00000003_sig000005c9
    );
  blk00000003_blk0000037e : XORCY
    port map (
      CI => blk00000003_sig000005c4,
      LI => blk00000003_sig000005c5,
      O => blk00000003_sig000005c6
    );
  blk00000003_blk0000037d : XORCY
    port map (
      CI => blk00000003_sig000005c1,
      LI => blk00000003_sig000005c2,
      O => blk00000003_sig000005c3
    );
  blk00000003_blk0000037c : XORCY
    port map (
      CI => blk00000003_sig000005be,
      LI => blk00000003_sig000005bf,
      O => blk00000003_sig000005c0
    );
  blk00000003_blk0000037b : XORCY
    port map (
      CI => blk00000003_sig000005bb,
      LI => blk00000003_sig000005bc,
      O => blk00000003_sig000005bd
    );
  blk00000003_blk0000037a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005b6,
      Q => blk00000003_sig000005ba
    );
  blk00000003_blk00000379 : MUXCY
    port map (
      CI => blk00000003_sig000005b7,
      DI => blk00000003_sig00000048,
      S => blk00000003_sig000005b8,
      O => blk00000003_sig000005a3
    );
  blk00000003_blk00000378 : XORCY
    port map (
      CI => blk00000003_sig000005b7,
      LI => blk00000003_sig000005b8,
      O => blk00000003_sig000005b9
    );
  blk00000003_blk00000377 : MUXCY
    port map (
      CI => blk00000003_sig00000576,
      DI => blk00000003_sig000005b5,
      S => blk00000003_sig00000577,
      O => blk00000003_sig000005b6
    );
  blk00000003_blk00000376 : MUXCY
    port map (
      CI => blk00000003_sig000005a3,
      DI => blk00000003_sig000005b4,
      S => blk00000003_sig000005a4,
      O => blk00000003_sig000005a0
    );
  blk00000003_blk00000375 : MUXCY
    port map (
      CI => blk00000003_sig000005a0,
      DI => blk00000003_sig000005b3,
      S => blk00000003_sig000005a1,
      O => blk00000003_sig0000059d
    );
  blk00000003_blk00000374 : MUXCY
    port map (
      CI => blk00000003_sig0000059d,
      DI => blk00000003_sig000005b2,
      S => blk00000003_sig0000059e,
      O => blk00000003_sig0000059a
    );
  blk00000003_blk00000373 : MUXCY
    port map (
      CI => blk00000003_sig0000059a,
      DI => blk00000003_sig000005b1,
      S => blk00000003_sig0000059b,
      O => blk00000003_sig00000597
    );
  blk00000003_blk00000372 : MUXCY
    port map (
      CI => blk00000003_sig00000597,
      DI => blk00000003_sig000005b0,
      S => blk00000003_sig00000598,
      O => blk00000003_sig00000594
    );
  blk00000003_blk00000371 : MUXCY
    port map (
      CI => blk00000003_sig00000594,
      DI => blk00000003_sig000005af,
      S => blk00000003_sig00000595,
      O => blk00000003_sig00000591
    );
  blk00000003_blk00000370 : MUXCY
    port map (
      CI => blk00000003_sig00000591,
      DI => blk00000003_sig000005ae,
      S => blk00000003_sig00000592,
      O => blk00000003_sig0000058e
    );
  blk00000003_blk0000036f : MUXCY
    port map (
      CI => blk00000003_sig0000058e,
      DI => blk00000003_sig000005ad,
      S => blk00000003_sig0000058f,
      O => blk00000003_sig0000058b
    );
  blk00000003_blk0000036e : MUXCY
    port map (
      CI => blk00000003_sig0000058b,
      DI => blk00000003_sig000005ac,
      S => blk00000003_sig0000058c,
      O => blk00000003_sig00000588
    );
  blk00000003_blk0000036d : MUXCY
    port map (
      CI => blk00000003_sig00000588,
      DI => blk00000003_sig000005ab,
      S => blk00000003_sig00000589,
      O => blk00000003_sig00000585
    );
  blk00000003_blk0000036c : MUXCY
    port map (
      CI => blk00000003_sig00000585,
      DI => blk00000003_sig000005aa,
      S => blk00000003_sig00000586,
      O => blk00000003_sig00000582
    );
  blk00000003_blk0000036b : MUXCY
    port map (
      CI => blk00000003_sig00000582,
      DI => blk00000003_sig000005a9,
      S => blk00000003_sig00000583,
      O => blk00000003_sig0000057f
    );
  blk00000003_blk0000036a : MUXCY
    port map (
      CI => blk00000003_sig0000057f,
      DI => blk00000003_sig000005a8,
      S => blk00000003_sig00000580,
      O => blk00000003_sig0000057c
    );
  blk00000003_blk00000369 : MUXCY
    port map (
      CI => blk00000003_sig0000057c,
      DI => blk00000003_sig000005a7,
      S => blk00000003_sig0000057d,
      O => blk00000003_sig00000579
    );
  blk00000003_blk00000368 : MUXCY
    port map (
      CI => blk00000003_sig00000579,
      DI => blk00000003_sig000005a6,
      S => blk00000003_sig0000057a,
      O => blk00000003_sig00000576
    );
  blk00000003_blk00000367 : XORCY
    port map (
      CI => blk00000003_sig000005a3,
      LI => blk00000003_sig000005a4,
      O => blk00000003_sig000005a5
    );
  blk00000003_blk00000366 : XORCY
    port map (
      CI => blk00000003_sig000005a0,
      LI => blk00000003_sig000005a1,
      O => blk00000003_sig000005a2
    );
  blk00000003_blk00000365 : XORCY
    port map (
      CI => blk00000003_sig0000059d,
      LI => blk00000003_sig0000059e,
      O => blk00000003_sig0000059f
    );
  blk00000003_blk00000364 : XORCY
    port map (
      CI => blk00000003_sig0000059a,
      LI => blk00000003_sig0000059b,
      O => blk00000003_sig0000059c
    );
  blk00000003_blk00000363 : XORCY
    port map (
      CI => blk00000003_sig00000597,
      LI => blk00000003_sig00000598,
      O => blk00000003_sig00000599
    );
  blk00000003_blk00000362 : XORCY
    port map (
      CI => blk00000003_sig00000594,
      LI => blk00000003_sig00000595,
      O => blk00000003_sig00000596
    );
  blk00000003_blk00000361 : XORCY
    port map (
      CI => blk00000003_sig00000591,
      LI => blk00000003_sig00000592,
      O => blk00000003_sig00000593
    );
  blk00000003_blk00000360 : XORCY
    port map (
      CI => blk00000003_sig0000058e,
      LI => blk00000003_sig0000058f,
      O => blk00000003_sig00000590
    );
  blk00000003_blk0000035f : XORCY
    port map (
      CI => blk00000003_sig0000058b,
      LI => blk00000003_sig0000058c,
      O => blk00000003_sig0000058d
    );
  blk00000003_blk0000035e : XORCY
    port map (
      CI => blk00000003_sig00000588,
      LI => blk00000003_sig00000589,
      O => blk00000003_sig0000058a
    );
  blk00000003_blk0000035d : XORCY
    port map (
      CI => blk00000003_sig00000585,
      LI => blk00000003_sig00000586,
      O => blk00000003_sig00000587
    );
  blk00000003_blk0000035c : XORCY
    port map (
      CI => blk00000003_sig00000582,
      LI => blk00000003_sig00000583,
      O => blk00000003_sig00000584
    );
  blk00000003_blk0000035b : XORCY
    port map (
      CI => blk00000003_sig0000057f,
      LI => blk00000003_sig00000580,
      O => blk00000003_sig00000581
    );
  blk00000003_blk0000035a : XORCY
    port map (
      CI => blk00000003_sig0000057c,
      LI => blk00000003_sig0000057d,
      O => blk00000003_sig0000057e
    );
  blk00000003_blk00000359 : XORCY
    port map (
      CI => blk00000003_sig00000579,
      LI => blk00000003_sig0000057a,
      O => blk00000003_sig0000057b
    );
  blk00000003_blk00000358 : XORCY
    port map (
      CI => blk00000003_sig00000576,
      LI => blk00000003_sig00000577,
      O => blk00000003_sig00000578
    );
  blk00000003_blk00000357 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000571,
      Q => blk00000003_sig00000575
    );
  blk00000003_blk00000356 : MUXCY
    port map (
      CI => blk00000003_sig00000572,
      DI => blk00000003_sig0000004c,
      S => blk00000003_sig00000573,
      O => blk00000003_sig0000055e
    );
  blk00000003_blk00000355 : XORCY
    port map (
      CI => blk00000003_sig00000572,
      LI => blk00000003_sig00000573,
      O => blk00000003_sig00000574
    );
  blk00000003_blk00000354 : MUXCY
    port map (
      CI => blk00000003_sig00000531,
      DI => blk00000003_sig00000570,
      S => blk00000003_sig00000532,
      O => blk00000003_sig00000571
    );
  blk00000003_blk00000353 : MUXCY
    port map (
      CI => blk00000003_sig0000055e,
      DI => blk00000003_sig0000056f,
      S => blk00000003_sig0000055f,
      O => blk00000003_sig0000055b
    );
  blk00000003_blk00000352 : MUXCY
    port map (
      CI => blk00000003_sig0000055b,
      DI => blk00000003_sig0000056e,
      S => blk00000003_sig0000055c,
      O => blk00000003_sig00000558
    );
  blk00000003_blk00000351 : MUXCY
    port map (
      CI => blk00000003_sig00000558,
      DI => blk00000003_sig0000056d,
      S => blk00000003_sig00000559,
      O => blk00000003_sig00000555
    );
  blk00000003_blk00000350 : MUXCY
    port map (
      CI => blk00000003_sig00000555,
      DI => blk00000003_sig0000056c,
      S => blk00000003_sig00000556,
      O => blk00000003_sig00000552
    );
  blk00000003_blk0000034f : MUXCY
    port map (
      CI => blk00000003_sig00000552,
      DI => blk00000003_sig0000056b,
      S => blk00000003_sig00000553,
      O => blk00000003_sig0000054f
    );
  blk00000003_blk0000034e : MUXCY
    port map (
      CI => blk00000003_sig0000054f,
      DI => blk00000003_sig0000056a,
      S => blk00000003_sig00000550,
      O => blk00000003_sig0000054c
    );
  blk00000003_blk0000034d : MUXCY
    port map (
      CI => blk00000003_sig0000054c,
      DI => blk00000003_sig00000569,
      S => blk00000003_sig0000054d,
      O => blk00000003_sig00000549
    );
  blk00000003_blk0000034c : MUXCY
    port map (
      CI => blk00000003_sig00000549,
      DI => blk00000003_sig00000568,
      S => blk00000003_sig0000054a,
      O => blk00000003_sig00000546
    );
  blk00000003_blk0000034b : MUXCY
    port map (
      CI => blk00000003_sig00000546,
      DI => blk00000003_sig00000567,
      S => blk00000003_sig00000547,
      O => blk00000003_sig00000543
    );
  blk00000003_blk0000034a : MUXCY
    port map (
      CI => blk00000003_sig00000543,
      DI => blk00000003_sig00000566,
      S => blk00000003_sig00000544,
      O => blk00000003_sig00000540
    );
  blk00000003_blk00000349 : MUXCY
    port map (
      CI => blk00000003_sig00000540,
      DI => blk00000003_sig00000565,
      S => blk00000003_sig00000541,
      O => blk00000003_sig0000053d
    );
  blk00000003_blk00000348 : MUXCY
    port map (
      CI => blk00000003_sig0000053d,
      DI => blk00000003_sig00000564,
      S => blk00000003_sig0000053e,
      O => blk00000003_sig0000053a
    );
  blk00000003_blk00000347 : MUXCY
    port map (
      CI => blk00000003_sig0000053a,
      DI => blk00000003_sig00000563,
      S => blk00000003_sig0000053b,
      O => blk00000003_sig00000537
    );
  blk00000003_blk00000346 : MUXCY
    port map (
      CI => blk00000003_sig00000537,
      DI => blk00000003_sig00000562,
      S => blk00000003_sig00000538,
      O => blk00000003_sig00000534
    );
  blk00000003_blk00000345 : MUXCY
    port map (
      CI => blk00000003_sig00000534,
      DI => blk00000003_sig00000561,
      S => blk00000003_sig00000535,
      O => blk00000003_sig00000531
    );
  blk00000003_blk00000344 : XORCY
    port map (
      CI => blk00000003_sig0000055e,
      LI => blk00000003_sig0000055f,
      O => blk00000003_sig00000560
    );
  blk00000003_blk00000343 : XORCY
    port map (
      CI => blk00000003_sig0000055b,
      LI => blk00000003_sig0000055c,
      O => blk00000003_sig0000055d
    );
  blk00000003_blk00000342 : XORCY
    port map (
      CI => blk00000003_sig00000558,
      LI => blk00000003_sig00000559,
      O => blk00000003_sig0000055a
    );
  blk00000003_blk00000341 : XORCY
    port map (
      CI => blk00000003_sig00000555,
      LI => blk00000003_sig00000556,
      O => blk00000003_sig00000557
    );
  blk00000003_blk00000340 : XORCY
    port map (
      CI => blk00000003_sig00000552,
      LI => blk00000003_sig00000553,
      O => blk00000003_sig00000554
    );
  blk00000003_blk0000033f : XORCY
    port map (
      CI => blk00000003_sig0000054f,
      LI => blk00000003_sig00000550,
      O => blk00000003_sig00000551
    );
  blk00000003_blk0000033e : XORCY
    port map (
      CI => blk00000003_sig0000054c,
      LI => blk00000003_sig0000054d,
      O => blk00000003_sig0000054e
    );
  blk00000003_blk0000033d : XORCY
    port map (
      CI => blk00000003_sig00000549,
      LI => blk00000003_sig0000054a,
      O => blk00000003_sig0000054b
    );
  blk00000003_blk0000033c : XORCY
    port map (
      CI => blk00000003_sig00000546,
      LI => blk00000003_sig00000547,
      O => blk00000003_sig00000548
    );
  blk00000003_blk0000033b : XORCY
    port map (
      CI => blk00000003_sig00000543,
      LI => blk00000003_sig00000544,
      O => blk00000003_sig00000545
    );
  blk00000003_blk0000033a : XORCY
    port map (
      CI => blk00000003_sig00000540,
      LI => blk00000003_sig00000541,
      O => blk00000003_sig00000542
    );
  blk00000003_blk00000339 : XORCY
    port map (
      CI => blk00000003_sig0000053d,
      LI => blk00000003_sig0000053e,
      O => blk00000003_sig0000053f
    );
  blk00000003_blk00000338 : XORCY
    port map (
      CI => blk00000003_sig0000053a,
      LI => blk00000003_sig0000053b,
      O => blk00000003_sig0000053c
    );
  blk00000003_blk00000337 : XORCY
    port map (
      CI => blk00000003_sig00000537,
      LI => blk00000003_sig00000538,
      O => blk00000003_sig00000539
    );
  blk00000003_blk00000336 : XORCY
    port map (
      CI => blk00000003_sig00000534,
      LI => blk00000003_sig00000535,
      O => blk00000003_sig00000536
    );
  blk00000003_blk00000335 : XORCY
    port map (
      CI => blk00000003_sig00000531,
      LI => blk00000003_sig00000532,
      O => blk00000003_sig00000533
    );
  blk00000003_blk00000334 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000052c,
      Q => blk00000003_sig00000530
    );
  blk00000003_blk00000333 : MUXCY
    port map (
      CI => blk00000003_sig0000052d,
      DI => blk00000003_sig00000051,
      S => blk00000003_sig0000052e,
      O => blk00000003_sig00000519
    );
  blk00000003_blk00000332 : XORCY
    port map (
      CI => blk00000003_sig0000052d,
      LI => blk00000003_sig0000052e,
      O => blk00000003_sig0000052f
    );
  blk00000003_blk00000331 : MUXCY
    port map (
      CI => blk00000003_sig000004ec,
      DI => blk00000003_sig0000052b,
      S => blk00000003_sig000004ed,
      O => blk00000003_sig0000052c
    );
  blk00000003_blk00000330 : MUXCY
    port map (
      CI => blk00000003_sig00000519,
      DI => blk00000003_sig0000052a,
      S => blk00000003_sig0000051a,
      O => blk00000003_sig00000516
    );
  blk00000003_blk0000032f : MUXCY
    port map (
      CI => blk00000003_sig00000516,
      DI => blk00000003_sig00000529,
      S => blk00000003_sig00000517,
      O => blk00000003_sig00000513
    );
  blk00000003_blk0000032e : MUXCY
    port map (
      CI => blk00000003_sig00000513,
      DI => blk00000003_sig00000528,
      S => blk00000003_sig00000514,
      O => blk00000003_sig00000510
    );
  blk00000003_blk0000032d : MUXCY
    port map (
      CI => blk00000003_sig00000510,
      DI => blk00000003_sig00000527,
      S => blk00000003_sig00000511,
      O => blk00000003_sig0000050d
    );
  blk00000003_blk0000032c : MUXCY
    port map (
      CI => blk00000003_sig0000050d,
      DI => blk00000003_sig00000526,
      S => blk00000003_sig0000050e,
      O => blk00000003_sig0000050a
    );
  blk00000003_blk0000032b : MUXCY
    port map (
      CI => blk00000003_sig0000050a,
      DI => blk00000003_sig00000525,
      S => blk00000003_sig0000050b,
      O => blk00000003_sig00000507
    );
  blk00000003_blk0000032a : MUXCY
    port map (
      CI => blk00000003_sig00000507,
      DI => blk00000003_sig00000524,
      S => blk00000003_sig00000508,
      O => blk00000003_sig00000504
    );
  blk00000003_blk00000329 : MUXCY
    port map (
      CI => blk00000003_sig00000504,
      DI => blk00000003_sig00000523,
      S => blk00000003_sig00000505,
      O => blk00000003_sig00000501
    );
  blk00000003_blk00000328 : MUXCY
    port map (
      CI => blk00000003_sig00000501,
      DI => blk00000003_sig00000522,
      S => blk00000003_sig00000502,
      O => blk00000003_sig000004fe
    );
  blk00000003_blk00000327 : MUXCY
    port map (
      CI => blk00000003_sig000004fe,
      DI => blk00000003_sig00000521,
      S => blk00000003_sig000004ff,
      O => blk00000003_sig000004fb
    );
  blk00000003_blk00000326 : MUXCY
    port map (
      CI => blk00000003_sig000004fb,
      DI => blk00000003_sig00000520,
      S => blk00000003_sig000004fc,
      O => blk00000003_sig000004f8
    );
  blk00000003_blk00000325 : MUXCY
    port map (
      CI => blk00000003_sig000004f8,
      DI => blk00000003_sig0000051f,
      S => blk00000003_sig000004f9,
      O => blk00000003_sig000004f5
    );
  blk00000003_blk00000324 : MUXCY
    port map (
      CI => blk00000003_sig000004f5,
      DI => blk00000003_sig0000051e,
      S => blk00000003_sig000004f6,
      O => blk00000003_sig000004f2
    );
  blk00000003_blk00000323 : MUXCY
    port map (
      CI => blk00000003_sig000004f2,
      DI => blk00000003_sig0000051d,
      S => blk00000003_sig000004f3,
      O => blk00000003_sig000004ef
    );
  blk00000003_blk00000322 : MUXCY
    port map (
      CI => blk00000003_sig000004ef,
      DI => blk00000003_sig0000051c,
      S => blk00000003_sig000004f0,
      O => blk00000003_sig000004ec
    );
  blk00000003_blk00000321 : XORCY
    port map (
      CI => blk00000003_sig00000519,
      LI => blk00000003_sig0000051a,
      O => blk00000003_sig0000051b
    );
  blk00000003_blk00000320 : XORCY
    port map (
      CI => blk00000003_sig00000516,
      LI => blk00000003_sig00000517,
      O => blk00000003_sig00000518
    );
  blk00000003_blk0000031f : XORCY
    port map (
      CI => blk00000003_sig00000513,
      LI => blk00000003_sig00000514,
      O => blk00000003_sig00000515
    );
  blk00000003_blk0000031e : XORCY
    port map (
      CI => blk00000003_sig00000510,
      LI => blk00000003_sig00000511,
      O => blk00000003_sig00000512
    );
  blk00000003_blk0000031d : XORCY
    port map (
      CI => blk00000003_sig0000050d,
      LI => blk00000003_sig0000050e,
      O => blk00000003_sig0000050f
    );
  blk00000003_blk0000031c : XORCY
    port map (
      CI => blk00000003_sig0000050a,
      LI => blk00000003_sig0000050b,
      O => blk00000003_sig0000050c
    );
  blk00000003_blk0000031b : XORCY
    port map (
      CI => blk00000003_sig00000507,
      LI => blk00000003_sig00000508,
      O => blk00000003_sig00000509
    );
  blk00000003_blk0000031a : XORCY
    port map (
      CI => blk00000003_sig00000504,
      LI => blk00000003_sig00000505,
      O => blk00000003_sig00000506
    );
  blk00000003_blk00000319 : XORCY
    port map (
      CI => blk00000003_sig00000501,
      LI => blk00000003_sig00000502,
      O => blk00000003_sig00000503
    );
  blk00000003_blk00000318 : XORCY
    port map (
      CI => blk00000003_sig000004fe,
      LI => blk00000003_sig000004ff,
      O => blk00000003_sig00000500
    );
  blk00000003_blk00000317 : XORCY
    port map (
      CI => blk00000003_sig000004fb,
      LI => blk00000003_sig000004fc,
      O => blk00000003_sig000004fd
    );
  blk00000003_blk00000316 : XORCY
    port map (
      CI => blk00000003_sig000004f8,
      LI => blk00000003_sig000004f9,
      O => blk00000003_sig000004fa
    );
  blk00000003_blk00000315 : XORCY
    port map (
      CI => blk00000003_sig000004f5,
      LI => blk00000003_sig000004f6,
      O => blk00000003_sig000004f7
    );
  blk00000003_blk00000314 : XORCY
    port map (
      CI => blk00000003_sig000004f2,
      LI => blk00000003_sig000004f3,
      O => blk00000003_sig000004f4
    );
  blk00000003_blk00000313 : XORCY
    port map (
      CI => blk00000003_sig000004ef,
      LI => blk00000003_sig000004f0,
      O => blk00000003_sig000004f1
    );
  blk00000003_blk00000312 : XORCY
    port map (
      CI => blk00000003_sig000004ec,
      LI => blk00000003_sig000004ed,
      O => blk00000003_sig000004ee
    );
  blk00000003_blk00000311 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004e7,
      Q => blk00000003_sig000004eb
    );
  blk00000003_blk00000310 : MUXCY
    port map (
      CI => blk00000003_sig000004e8,
      DI => blk00000003_sig00000057,
      S => blk00000003_sig000004e9,
      O => blk00000003_sig000004d4
    );
  blk00000003_blk0000030f : XORCY
    port map (
      CI => blk00000003_sig000004e8,
      LI => blk00000003_sig000004e9,
      O => blk00000003_sig000004ea
    );
  blk00000003_blk0000030e : MUXCY
    port map (
      CI => blk00000003_sig000004a7,
      DI => blk00000003_sig000004e6,
      S => blk00000003_sig000004a8,
      O => blk00000003_sig000004e7
    );
  blk00000003_blk0000030d : MUXCY
    port map (
      CI => blk00000003_sig000004d4,
      DI => blk00000003_sig000004e5,
      S => blk00000003_sig000004d5,
      O => blk00000003_sig000004d1
    );
  blk00000003_blk0000030c : MUXCY
    port map (
      CI => blk00000003_sig000004d1,
      DI => blk00000003_sig000004e4,
      S => blk00000003_sig000004d2,
      O => blk00000003_sig000004ce
    );
  blk00000003_blk0000030b : MUXCY
    port map (
      CI => blk00000003_sig000004ce,
      DI => blk00000003_sig000004e3,
      S => blk00000003_sig000004cf,
      O => blk00000003_sig000004cb
    );
  blk00000003_blk0000030a : MUXCY
    port map (
      CI => blk00000003_sig000004cb,
      DI => blk00000003_sig000004e2,
      S => blk00000003_sig000004cc,
      O => blk00000003_sig000004c8
    );
  blk00000003_blk00000309 : MUXCY
    port map (
      CI => blk00000003_sig000004c8,
      DI => blk00000003_sig000004e1,
      S => blk00000003_sig000004c9,
      O => blk00000003_sig000004c5
    );
  blk00000003_blk00000308 : MUXCY
    port map (
      CI => blk00000003_sig000004c5,
      DI => blk00000003_sig000004e0,
      S => blk00000003_sig000004c6,
      O => blk00000003_sig000004c2
    );
  blk00000003_blk00000307 : MUXCY
    port map (
      CI => blk00000003_sig000004c2,
      DI => blk00000003_sig000004df,
      S => blk00000003_sig000004c3,
      O => blk00000003_sig000004bf
    );
  blk00000003_blk00000306 : MUXCY
    port map (
      CI => blk00000003_sig000004bf,
      DI => blk00000003_sig000004de,
      S => blk00000003_sig000004c0,
      O => blk00000003_sig000004bc
    );
  blk00000003_blk00000305 : MUXCY
    port map (
      CI => blk00000003_sig000004bc,
      DI => blk00000003_sig000004dd,
      S => blk00000003_sig000004bd,
      O => blk00000003_sig000004b9
    );
  blk00000003_blk00000304 : MUXCY
    port map (
      CI => blk00000003_sig000004b9,
      DI => blk00000003_sig000004dc,
      S => blk00000003_sig000004ba,
      O => blk00000003_sig000004b6
    );
  blk00000003_blk00000303 : MUXCY
    port map (
      CI => blk00000003_sig000004b6,
      DI => blk00000003_sig000004db,
      S => blk00000003_sig000004b7,
      O => blk00000003_sig000004b3
    );
  blk00000003_blk00000302 : MUXCY
    port map (
      CI => blk00000003_sig000004b3,
      DI => blk00000003_sig000004da,
      S => blk00000003_sig000004b4,
      O => blk00000003_sig000004b0
    );
  blk00000003_blk00000301 : MUXCY
    port map (
      CI => blk00000003_sig000004b0,
      DI => blk00000003_sig000004d9,
      S => blk00000003_sig000004b1,
      O => blk00000003_sig000004ad
    );
  blk00000003_blk00000300 : MUXCY
    port map (
      CI => blk00000003_sig000004ad,
      DI => blk00000003_sig000004d8,
      S => blk00000003_sig000004ae,
      O => blk00000003_sig000004aa
    );
  blk00000003_blk000002ff : MUXCY
    port map (
      CI => blk00000003_sig000004aa,
      DI => blk00000003_sig000004d7,
      S => blk00000003_sig000004ab,
      O => blk00000003_sig000004a7
    );
  blk00000003_blk000002fe : XORCY
    port map (
      CI => blk00000003_sig000004d4,
      LI => blk00000003_sig000004d5,
      O => blk00000003_sig000004d6
    );
  blk00000003_blk000002fd : XORCY
    port map (
      CI => blk00000003_sig000004d1,
      LI => blk00000003_sig000004d2,
      O => blk00000003_sig000004d3
    );
  blk00000003_blk000002fc : XORCY
    port map (
      CI => blk00000003_sig000004ce,
      LI => blk00000003_sig000004cf,
      O => blk00000003_sig000004d0
    );
  blk00000003_blk000002fb : XORCY
    port map (
      CI => blk00000003_sig000004cb,
      LI => blk00000003_sig000004cc,
      O => blk00000003_sig000004cd
    );
  blk00000003_blk000002fa : XORCY
    port map (
      CI => blk00000003_sig000004c8,
      LI => blk00000003_sig000004c9,
      O => blk00000003_sig000004ca
    );
  blk00000003_blk000002f9 : XORCY
    port map (
      CI => blk00000003_sig000004c5,
      LI => blk00000003_sig000004c6,
      O => blk00000003_sig000004c7
    );
  blk00000003_blk000002f8 : XORCY
    port map (
      CI => blk00000003_sig000004c2,
      LI => blk00000003_sig000004c3,
      O => blk00000003_sig000004c4
    );
  blk00000003_blk000002f7 : XORCY
    port map (
      CI => blk00000003_sig000004bf,
      LI => blk00000003_sig000004c0,
      O => blk00000003_sig000004c1
    );
  blk00000003_blk000002f6 : XORCY
    port map (
      CI => blk00000003_sig000004bc,
      LI => blk00000003_sig000004bd,
      O => blk00000003_sig000004be
    );
  blk00000003_blk000002f5 : XORCY
    port map (
      CI => blk00000003_sig000004b9,
      LI => blk00000003_sig000004ba,
      O => blk00000003_sig000004bb
    );
  blk00000003_blk000002f4 : XORCY
    port map (
      CI => blk00000003_sig000004b6,
      LI => blk00000003_sig000004b7,
      O => blk00000003_sig000004b8
    );
  blk00000003_blk000002f3 : XORCY
    port map (
      CI => blk00000003_sig000004b3,
      LI => blk00000003_sig000004b4,
      O => blk00000003_sig000004b5
    );
  blk00000003_blk000002f2 : XORCY
    port map (
      CI => blk00000003_sig000004b0,
      LI => blk00000003_sig000004b1,
      O => blk00000003_sig000004b2
    );
  blk00000003_blk000002f1 : XORCY
    port map (
      CI => blk00000003_sig000004ad,
      LI => blk00000003_sig000004ae,
      O => blk00000003_sig000004af
    );
  blk00000003_blk000002f0 : XORCY
    port map (
      CI => blk00000003_sig000004aa,
      LI => blk00000003_sig000004ab,
      O => blk00000003_sig000004ac
    );
  blk00000003_blk000002ef : XORCY
    port map (
      CI => blk00000003_sig000004a7,
      LI => blk00000003_sig000004a8,
      O => blk00000003_sig000004a9
    );
  blk00000003_blk000002ee : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004a2,
      Q => blk00000003_sig000004a6
    );
  blk00000003_blk000002ed : MUXCY
    port map (
      CI => blk00000003_sig000004a3,
      DI => blk00000003_sig0000005e,
      S => blk00000003_sig000004a4,
      O => blk00000003_sig0000048f
    );
  blk00000003_blk000002ec : XORCY
    port map (
      CI => blk00000003_sig000004a3,
      LI => blk00000003_sig000004a4,
      O => blk00000003_sig000004a5
    );
  blk00000003_blk000002eb : MUXCY
    port map (
      CI => blk00000003_sig00000462,
      DI => blk00000003_sig000004a1,
      S => blk00000003_sig00000463,
      O => blk00000003_sig000004a2
    );
  blk00000003_blk000002ea : MUXCY
    port map (
      CI => blk00000003_sig0000048f,
      DI => blk00000003_sig000004a0,
      S => blk00000003_sig00000490,
      O => blk00000003_sig0000048c
    );
  blk00000003_blk000002e9 : MUXCY
    port map (
      CI => blk00000003_sig0000048c,
      DI => blk00000003_sig0000049f,
      S => blk00000003_sig0000048d,
      O => blk00000003_sig00000489
    );
  blk00000003_blk000002e8 : MUXCY
    port map (
      CI => blk00000003_sig00000489,
      DI => blk00000003_sig0000049e,
      S => blk00000003_sig0000048a,
      O => blk00000003_sig00000486
    );
  blk00000003_blk000002e7 : MUXCY
    port map (
      CI => blk00000003_sig00000486,
      DI => blk00000003_sig0000049d,
      S => blk00000003_sig00000487,
      O => blk00000003_sig00000483
    );
  blk00000003_blk000002e6 : MUXCY
    port map (
      CI => blk00000003_sig00000483,
      DI => blk00000003_sig0000049c,
      S => blk00000003_sig00000484,
      O => blk00000003_sig00000480
    );
  blk00000003_blk000002e5 : MUXCY
    port map (
      CI => blk00000003_sig00000480,
      DI => blk00000003_sig0000049b,
      S => blk00000003_sig00000481,
      O => blk00000003_sig0000047d
    );
  blk00000003_blk000002e4 : MUXCY
    port map (
      CI => blk00000003_sig0000047d,
      DI => blk00000003_sig0000049a,
      S => blk00000003_sig0000047e,
      O => blk00000003_sig0000047a
    );
  blk00000003_blk000002e3 : MUXCY
    port map (
      CI => blk00000003_sig0000047a,
      DI => blk00000003_sig00000499,
      S => blk00000003_sig0000047b,
      O => blk00000003_sig00000477
    );
  blk00000003_blk000002e2 : MUXCY
    port map (
      CI => blk00000003_sig00000477,
      DI => blk00000003_sig00000498,
      S => blk00000003_sig00000478,
      O => blk00000003_sig00000474
    );
  blk00000003_blk000002e1 : MUXCY
    port map (
      CI => blk00000003_sig00000474,
      DI => blk00000003_sig00000497,
      S => blk00000003_sig00000475,
      O => blk00000003_sig00000471
    );
  blk00000003_blk000002e0 : MUXCY
    port map (
      CI => blk00000003_sig00000471,
      DI => blk00000003_sig00000496,
      S => blk00000003_sig00000472,
      O => blk00000003_sig0000046e
    );
  blk00000003_blk000002df : MUXCY
    port map (
      CI => blk00000003_sig0000046e,
      DI => blk00000003_sig00000495,
      S => blk00000003_sig0000046f,
      O => blk00000003_sig0000046b
    );
  blk00000003_blk000002de : MUXCY
    port map (
      CI => blk00000003_sig0000046b,
      DI => blk00000003_sig00000494,
      S => blk00000003_sig0000046c,
      O => blk00000003_sig00000468
    );
  blk00000003_blk000002dd : MUXCY
    port map (
      CI => blk00000003_sig00000468,
      DI => blk00000003_sig00000493,
      S => blk00000003_sig00000469,
      O => blk00000003_sig00000465
    );
  blk00000003_blk000002dc : MUXCY
    port map (
      CI => blk00000003_sig00000465,
      DI => blk00000003_sig00000492,
      S => blk00000003_sig00000466,
      O => blk00000003_sig00000462
    );
  blk00000003_blk000002db : XORCY
    port map (
      CI => blk00000003_sig0000048f,
      LI => blk00000003_sig00000490,
      O => blk00000003_sig00000491
    );
  blk00000003_blk000002da : XORCY
    port map (
      CI => blk00000003_sig0000048c,
      LI => blk00000003_sig0000048d,
      O => blk00000003_sig0000048e
    );
  blk00000003_blk000002d9 : XORCY
    port map (
      CI => blk00000003_sig00000489,
      LI => blk00000003_sig0000048a,
      O => blk00000003_sig0000048b
    );
  blk00000003_blk000002d8 : XORCY
    port map (
      CI => blk00000003_sig00000486,
      LI => blk00000003_sig00000487,
      O => blk00000003_sig00000488
    );
  blk00000003_blk000002d7 : XORCY
    port map (
      CI => blk00000003_sig00000483,
      LI => blk00000003_sig00000484,
      O => blk00000003_sig00000485
    );
  blk00000003_blk000002d6 : XORCY
    port map (
      CI => blk00000003_sig00000480,
      LI => blk00000003_sig00000481,
      O => blk00000003_sig00000482
    );
  blk00000003_blk000002d5 : XORCY
    port map (
      CI => blk00000003_sig0000047d,
      LI => blk00000003_sig0000047e,
      O => blk00000003_sig0000047f
    );
  blk00000003_blk000002d4 : XORCY
    port map (
      CI => blk00000003_sig0000047a,
      LI => blk00000003_sig0000047b,
      O => blk00000003_sig0000047c
    );
  blk00000003_blk000002d3 : XORCY
    port map (
      CI => blk00000003_sig00000477,
      LI => blk00000003_sig00000478,
      O => blk00000003_sig00000479
    );
  blk00000003_blk000002d2 : XORCY
    port map (
      CI => blk00000003_sig00000474,
      LI => blk00000003_sig00000475,
      O => blk00000003_sig00000476
    );
  blk00000003_blk000002d1 : XORCY
    port map (
      CI => blk00000003_sig00000471,
      LI => blk00000003_sig00000472,
      O => blk00000003_sig00000473
    );
  blk00000003_blk000002d0 : XORCY
    port map (
      CI => blk00000003_sig0000046e,
      LI => blk00000003_sig0000046f,
      O => blk00000003_sig00000470
    );
  blk00000003_blk000002cf : XORCY
    port map (
      CI => blk00000003_sig0000046b,
      LI => blk00000003_sig0000046c,
      O => blk00000003_sig0000046d
    );
  blk00000003_blk000002ce : XORCY
    port map (
      CI => blk00000003_sig00000468,
      LI => blk00000003_sig00000469,
      O => blk00000003_sig0000046a
    );
  blk00000003_blk000002cd : XORCY
    port map (
      CI => blk00000003_sig00000465,
      LI => blk00000003_sig00000466,
      O => blk00000003_sig00000467
    );
  blk00000003_blk000002cc : XORCY
    port map (
      CI => blk00000003_sig00000462,
      LI => blk00000003_sig00000463,
      O => blk00000003_sig00000464
    );
  blk00000003_blk000002cb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000045d,
      Q => blk00000003_sig00000461
    );
  blk00000003_blk000002ca : MUXCY
    port map (
      CI => blk00000003_sig0000045e,
      DI => blk00000003_sig00000066,
      S => blk00000003_sig0000045f,
      O => blk00000003_sig0000044a
    );
  blk00000003_blk000002c9 : XORCY
    port map (
      CI => blk00000003_sig0000045e,
      LI => blk00000003_sig0000045f,
      O => blk00000003_sig00000460
    );
  blk00000003_blk000002c8 : MUXCY
    port map (
      CI => blk00000003_sig0000041d,
      DI => blk00000003_sig0000045c,
      S => blk00000003_sig0000041e,
      O => blk00000003_sig0000045d
    );
  blk00000003_blk000002c7 : MUXCY
    port map (
      CI => blk00000003_sig0000044a,
      DI => blk00000003_sig0000045b,
      S => blk00000003_sig0000044b,
      O => blk00000003_sig00000447
    );
  blk00000003_blk000002c6 : MUXCY
    port map (
      CI => blk00000003_sig00000447,
      DI => blk00000003_sig0000045a,
      S => blk00000003_sig00000448,
      O => blk00000003_sig00000444
    );
  blk00000003_blk000002c5 : MUXCY
    port map (
      CI => blk00000003_sig00000444,
      DI => blk00000003_sig00000459,
      S => blk00000003_sig00000445,
      O => blk00000003_sig00000441
    );
  blk00000003_blk000002c4 : MUXCY
    port map (
      CI => blk00000003_sig00000441,
      DI => blk00000003_sig00000458,
      S => blk00000003_sig00000442,
      O => blk00000003_sig0000043e
    );
  blk00000003_blk000002c3 : MUXCY
    port map (
      CI => blk00000003_sig0000043e,
      DI => blk00000003_sig00000457,
      S => blk00000003_sig0000043f,
      O => blk00000003_sig0000043b
    );
  blk00000003_blk000002c2 : MUXCY
    port map (
      CI => blk00000003_sig0000043b,
      DI => blk00000003_sig00000456,
      S => blk00000003_sig0000043c,
      O => blk00000003_sig00000438
    );
  blk00000003_blk000002c1 : MUXCY
    port map (
      CI => blk00000003_sig00000438,
      DI => blk00000003_sig00000455,
      S => blk00000003_sig00000439,
      O => blk00000003_sig00000435
    );
  blk00000003_blk000002c0 : MUXCY
    port map (
      CI => blk00000003_sig00000435,
      DI => blk00000003_sig00000454,
      S => blk00000003_sig00000436,
      O => blk00000003_sig00000432
    );
  blk00000003_blk000002bf : MUXCY
    port map (
      CI => blk00000003_sig00000432,
      DI => blk00000003_sig00000453,
      S => blk00000003_sig00000433,
      O => blk00000003_sig0000042f
    );
  blk00000003_blk000002be : MUXCY
    port map (
      CI => blk00000003_sig0000042f,
      DI => blk00000003_sig00000452,
      S => blk00000003_sig00000430,
      O => blk00000003_sig0000042c
    );
  blk00000003_blk000002bd : MUXCY
    port map (
      CI => blk00000003_sig0000042c,
      DI => blk00000003_sig00000451,
      S => blk00000003_sig0000042d,
      O => blk00000003_sig00000429
    );
  blk00000003_blk000002bc : MUXCY
    port map (
      CI => blk00000003_sig00000429,
      DI => blk00000003_sig00000450,
      S => blk00000003_sig0000042a,
      O => blk00000003_sig00000426
    );
  blk00000003_blk000002bb : MUXCY
    port map (
      CI => blk00000003_sig00000426,
      DI => blk00000003_sig0000044f,
      S => blk00000003_sig00000427,
      O => blk00000003_sig00000423
    );
  blk00000003_blk000002ba : MUXCY
    port map (
      CI => blk00000003_sig00000423,
      DI => blk00000003_sig0000044e,
      S => blk00000003_sig00000424,
      O => blk00000003_sig00000420
    );
  blk00000003_blk000002b9 : MUXCY
    port map (
      CI => blk00000003_sig00000420,
      DI => blk00000003_sig0000044d,
      S => blk00000003_sig00000421,
      O => blk00000003_sig0000041d
    );
  blk00000003_blk000002b8 : XORCY
    port map (
      CI => blk00000003_sig0000044a,
      LI => blk00000003_sig0000044b,
      O => blk00000003_sig0000044c
    );
  blk00000003_blk000002b7 : XORCY
    port map (
      CI => blk00000003_sig00000447,
      LI => blk00000003_sig00000448,
      O => blk00000003_sig00000449
    );
  blk00000003_blk000002b6 : XORCY
    port map (
      CI => blk00000003_sig00000444,
      LI => blk00000003_sig00000445,
      O => blk00000003_sig00000446
    );
  blk00000003_blk000002b5 : XORCY
    port map (
      CI => blk00000003_sig00000441,
      LI => blk00000003_sig00000442,
      O => blk00000003_sig00000443
    );
  blk00000003_blk000002b4 : XORCY
    port map (
      CI => blk00000003_sig0000043e,
      LI => blk00000003_sig0000043f,
      O => blk00000003_sig00000440
    );
  blk00000003_blk000002b3 : XORCY
    port map (
      CI => blk00000003_sig0000043b,
      LI => blk00000003_sig0000043c,
      O => blk00000003_sig0000043d
    );
  blk00000003_blk000002b2 : XORCY
    port map (
      CI => blk00000003_sig00000438,
      LI => blk00000003_sig00000439,
      O => blk00000003_sig0000043a
    );
  blk00000003_blk000002b1 : XORCY
    port map (
      CI => blk00000003_sig00000435,
      LI => blk00000003_sig00000436,
      O => blk00000003_sig00000437
    );
  blk00000003_blk000002b0 : XORCY
    port map (
      CI => blk00000003_sig00000432,
      LI => blk00000003_sig00000433,
      O => blk00000003_sig00000434
    );
  blk00000003_blk000002af : XORCY
    port map (
      CI => blk00000003_sig0000042f,
      LI => blk00000003_sig00000430,
      O => blk00000003_sig00000431
    );
  blk00000003_blk000002ae : XORCY
    port map (
      CI => blk00000003_sig0000042c,
      LI => blk00000003_sig0000042d,
      O => blk00000003_sig0000042e
    );
  blk00000003_blk000002ad : XORCY
    port map (
      CI => blk00000003_sig00000429,
      LI => blk00000003_sig0000042a,
      O => blk00000003_sig0000042b
    );
  blk00000003_blk000002ac : XORCY
    port map (
      CI => blk00000003_sig00000426,
      LI => blk00000003_sig00000427,
      O => blk00000003_sig00000428
    );
  blk00000003_blk000002ab : XORCY
    port map (
      CI => blk00000003_sig00000423,
      LI => blk00000003_sig00000424,
      O => blk00000003_sig00000425
    );
  blk00000003_blk000002aa : XORCY
    port map (
      CI => blk00000003_sig00000420,
      LI => blk00000003_sig00000421,
      O => blk00000003_sig00000422
    );
  blk00000003_blk000002a9 : XORCY
    port map (
      CI => blk00000003_sig0000041d,
      LI => blk00000003_sig0000041e,
      O => blk00000003_sig0000041f
    );
  blk00000003_blk000002a8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000417,
      Q => blk00000003_sig0000041c
    );
  blk00000003_blk000002a7 : MUXCY
    port map (
      CI => blk00000003_sig00000418,
      DI => blk00000003_sig0000041b,
      S => blk00000003_sig00000419,
      O => blk00000003_sig00000404
    );
  blk00000003_blk000002a6 : XORCY
    port map (
      CI => blk00000003_sig00000418,
      LI => blk00000003_sig00000419,
      O => blk00000003_sig0000041a
    );
  blk00000003_blk000002a5 : MUXCY
    port map (
      CI => blk00000003_sig000003d7,
      DI => blk00000003_sig00000416,
      S => blk00000003_sig000003d8,
      O => blk00000003_sig00000417
    );
  blk00000003_blk000002a4 : MUXCY
    port map (
      CI => blk00000003_sig00000404,
      DI => blk00000003_sig00000415,
      S => blk00000003_sig00000405,
      O => blk00000003_sig00000401
    );
  blk00000003_blk000002a3 : MUXCY
    port map (
      CI => blk00000003_sig00000401,
      DI => blk00000003_sig00000414,
      S => blk00000003_sig00000402,
      O => blk00000003_sig000003fe
    );
  blk00000003_blk000002a2 : MUXCY
    port map (
      CI => blk00000003_sig000003fe,
      DI => blk00000003_sig00000413,
      S => blk00000003_sig000003ff,
      O => blk00000003_sig000003fb
    );
  blk00000003_blk000002a1 : MUXCY
    port map (
      CI => blk00000003_sig000003fb,
      DI => blk00000003_sig00000412,
      S => blk00000003_sig000003fc,
      O => blk00000003_sig000003f8
    );
  blk00000003_blk000002a0 : MUXCY
    port map (
      CI => blk00000003_sig000003f8,
      DI => blk00000003_sig00000411,
      S => blk00000003_sig000003f9,
      O => blk00000003_sig000003f5
    );
  blk00000003_blk0000029f : MUXCY
    port map (
      CI => blk00000003_sig000003f5,
      DI => blk00000003_sig00000410,
      S => blk00000003_sig000003f6,
      O => blk00000003_sig000003f2
    );
  blk00000003_blk0000029e : MUXCY
    port map (
      CI => blk00000003_sig000003f2,
      DI => blk00000003_sig0000040f,
      S => blk00000003_sig000003f3,
      O => blk00000003_sig000003ef
    );
  blk00000003_blk0000029d : MUXCY
    port map (
      CI => blk00000003_sig000003ef,
      DI => blk00000003_sig0000040e,
      S => blk00000003_sig000003f0,
      O => blk00000003_sig000003ec
    );
  blk00000003_blk0000029c : MUXCY
    port map (
      CI => blk00000003_sig000003ec,
      DI => blk00000003_sig0000040d,
      S => blk00000003_sig000003ed,
      O => blk00000003_sig000003e9
    );
  blk00000003_blk0000029b : MUXCY
    port map (
      CI => blk00000003_sig000003e9,
      DI => blk00000003_sig0000040c,
      S => blk00000003_sig000003ea,
      O => blk00000003_sig000003e6
    );
  blk00000003_blk0000029a : MUXCY
    port map (
      CI => blk00000003_sig000003e6,
      DI => blk00000003_sig0000040b,
      S => blk00000003_sig000003e7,
      O => blk00000003_sig000003e3
    );
  blk00000003_blk00000299 : MUXCY
    port map (
      CI => blk00000003_sig000003e3,
      DI => blk00000003_sig0000040a,
      S => blk00000003_sig000003e4,
      O => blk00000003_sig000003e0
    );
  blk00000003_blk00000298 : MUXCY
    port map (
      CI => blk00000003_sig000003e0,
      DI => blk00000003_sig00000409,
      S => blk00000003_sig000003e1,
      O => blk00000003_sig000003dd
    );
  blk00000003_blk00000297 : MUXCY
    port map (
      CI => blk00000003_sig000003dd,
      DI => blk00000003_sig00000408,
      S => blk00000003_sig000003de,
      O => blk00000003_sig000003da
    );
  blk00000003_blk00000296 : MUXCY
    port map (
      CI => blk00000003_sig000003da,
      DI => blk00000003_sig00000407,
      S => blk00000003_sig000003db,
      O => blk00000003_sig000003d7
    );
  blk00000003_blk00000295 : XORCY
    port map (
      CI => blk00000003_sig00000404,
      LI => blk00000003_sig00000405,
      O => blk00000003_sig00000406
    );
  blk00000003_blk00000294 : XORCY
    port map (
      CI => blk00000003_sig00000401,
      LI => blk00000003_sig00000402,
      O => blk00000003_sig00000403
    );
  blk00000003_blk00000293 : XORCY
    port map (
      CI => blk00000003_sig000003fe,
      LI => blk00000003_sig000003ff,
      O => blk00000003_sig00000400
    );
  blk00000003_blk00000292 : XORCY
    port map (
      CI => blk00000003_sig000003fb,
      LI => blk00000003_sig000003fc,
      O => blk00000003_sig000003fd
    );
  blk00000003_blk00000291 : XORCY
    port map (
      CI => blk00000003_sig000003f8,
      LI => blk00000003_sig000003f9,
      O => blk00000003_sig000003fa
    );
  blk00000003_blk00000290 : XORCY
    port map (
      CI => blk00000003_sig000003f5,
      LI => blk00000003_sig000003f6,
      O => blk00000003_sig000003f7
    );
  blk00000003_blk0000028f : XORCY
    port map (
      CI => blk00000003_sig000003f2,
      LI => blk00000003_sig000003f3,
      O => blk00000003_sig000003f4
    );
  blk00000003_blk0000028e : XORCY
    port map (
      CI => blk00000003_sig000003ef,
      LI => blk00000003_sig000003f0,
      O => blk00000003_sig000003f1
    );
  blk00000003_blk0000028d : XORCY
    port map (
      CI => blk00000003_sig000003ec,
      LI => blk00000003_sig000003ed,
      O => blk00000003_sig000003ee
    );
  blk00000003_blk0000028c : XORCY
    port map (
      CI => blk00000003_sig000003e9,
      LI => blk00000003_sig000003ea,
      O => blk00000003_sig000003eb
    );
  blk00000003_blk0000028b : XORCY
    port map (
      CI => blk00000003_sig000003e6,
      LI => blk00000003_sig000003e7,
      O => blk00000003_sig000003e8
    );
  blk00000003_blk0000028a : XORCY
    port map (
      CI => blk00000003_sig000003e3,
      LI => blk00000003_sig000003e4,
      O => blk00000003_sig000003e5
    );
  blk00000003_blk00000289 : XORCY
    port map (
      CI => blk00000003_sig000003e0,
      LI => blk00000003_sig000003e1,
      O => blk00000003_sig000003e2
    );
  blk00000003_blk00000288 : XORCY
    port map (
      CI => blk00000003_sig000003dd,
      LI => blk00000003_sig000003de,
      O => blk00000003_sig000003df
    );
  blk00000003_blk00000287 : XORCY
    port map (
      CI => blk00000003_sig000003da,
      LI => blk00000003_sig000003db,
      O => blk00000003_sig000003dc
    );
  blk00000003_blk00000286 : XORCY
    port map (
      CI => blk00000003_sig000003d7,
      LI => blk00000003_sig000003d8,
      O => blk00000003_sig000003d9
    );
  blk00000003_blk00000285 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003d1,
      Q => blk00000003_sig000003d6
    );
  blk00000003_blk00000284 : MUXCY
    port map (
      CI => blk00000003_sig000003d2,
      DI => blk00000003_sig000003d5,
      S => blk00000003_sig000003d3,
      O => blk00000003_sig000003be
    );
  blk00000003_blk00000283 : XORCY
    port map (
      CI => blk00000003_sig000003d2,
      LI => blk00000003_sig000003d3,
      O => blk00000003_sig000003d4
    );
  blk00000003_blk00000282 : MUXCY
    port map (
      CI => blk00000003_sig00000391,
      DI => blk00000003_sig000003d0,
      S => blk00000003_sig00000392,
      O => blk00000003_sig000003d1
    );
  blk00000003_blk00000281 : MUXCY
    port map (
      CI => blk00000003_sig000003be,
      DI => blk00000003_sig000003cf,
      S => blk00000003_sig000003bf,
      O => blk00000003_sig000003bb
    );
  blk00000003_blk00000280 : MUXCY
    port map (
      CI => blk00000003_sig000003bb,
      DI => blk00000003_sig000003ce,
      S => blk00000003_sig000003bc,
      O => blk00000003_sig000003b8
    );
  blk00000003_blk0000027f : MUXCY
    port map (
      CI => blk00000003_sig000003b8,
      DI => blk00000003_sig000003cd,
      S => blk00000003_sig000003b9,
      O => blk00000003_sig000003b5
    );
  blk00000003_blk0000027e : MUXCY
    port map (
      CI => blk00000003_sig000003b5,
      DI => blk00000003_sig000003cc,
      S => blk00000003_sig000003b6,
      O => blk00000003_sig000003b2
    );
  blk00000003_blk0000027d : MUXCY
    port map (
      CI => blk00000003_sig000003b2,
      DI => blk00000003_sig000003cb,
      S => blk00000003_sig000003b3,
      O => blk00000003_sig000003af
    );
  blk00000003_blk0000027c : MUXCY
    port map (
      CI => blk00000003_sig000003af,
      DI => blk00000003_sig000003ca,
      S => blk00000003_sig000003b0,
      O => blk00000003_sig000003ac
    );
  blk00000003_blk0000027b : MUXCY
    port map (
      CI => blk00000003_sig000003ac,
      DI => blk00000003_sig000003c9,
      S => blk00000003_sig000003ad,
      O => blk00000003_sig000003a9
    );
  blk00000003_blk0000027a : MUXCY
    port map (
      CI => blk00000003_sig000003a9,
      DI => blk00000003_sig000003c8,
      S => blk00000003_sig000003aa,
      O => blk00000003_sig000003a6
    );
  blk00000003_blk00000279 : MUXCY
    port map (
      CI => blk00000003_sig000003a6,
      DI => blk00000003_sig000003c7,
      S => blk00000003_sig000003a7,
      O => blk00000003_sig000003a3
    );
  blk00000003_blk00000278 : MUXCY
    port map (
      CI => blk00000003_sig000003a3,
      DI => blk00000003_sig000003c6,
      S => blk00000003_sig000003a4,
      O => blk00000003_sig000003a0
    );
  blk00000003_blk00000277 : MUXCY
    port map (
      CI => blk00000003_sig000003a0,
      DI => blk00000003_sig000003c5,
      S => blk00000003_sig000003a1,
      O => blk00000003_sig0000039d
    );
  blk00000003_blk00000276 : MUXCY
    port map (
      CI => blk00000003_sig0000039d,
      DI => blk00000003_sig000003c4,
      S => blk00000003_sig0000039e,
      O => blk00000003_sig0000039a
    );
  blk00000003_blk00000275 : MUXCY
    port map (
      CI => blk00000003_sig0000039a,
      DI => blk00000003_sig000003c3,
      S => blk00000003_sig0000039b,
      O => blk00000003_sig00000397
    );
  blk00000003_blk00000274 : MUXCY
    port map (
      CI => blk00000003_sig00000397,
      DI => blk00000003_sig000003c2,
      S => blk00000003_sig00000398,
      O => blk00000003_sig00000394
    );
  blk00000003_blk00000273 : MUXCY
    port map (
      CI => blk00000003_sig00000394,
      DI => blk00000003_sig000003c1,
      S => blk00000003_sig00000395,
      O => blk00000003_sig00000391
    );
  blk00000003_blk00000272 : XORCY
    port map (
      CI => blk00000003_sig000003be,
      LI => blk00000003_sig000003bf,
      O => blk00000003_sig000003c0
    );
  blk00000003_blk00000271 : XORCY
    port map (
      CI => blk00000003_sig000003bb,
      LI => blk00000003_sig000003bc,
      O => blk00000003_sig000003bd
    );
  blk00000003_blk00000270 : XORCY
    port map (
      CI => blk00000003_sig000003b8,
      LI => blk00000003_sig000003b9,
      O => blk00000003_sig000003ba
    );
  blk00000003_blk0000026f : XORCY
    port map (
      CI => blk00000003_sig000003b5,
      LI => blk00000003_sig000003b6,
      O => blk00000003_sig000003b7
    );
  blk00000003_blk0000026e : XORCY
    port map (
      CI => blk00000003_sig000003b2,
      LI => blk00000003_sig000003b3,
      O => blk00000003_sig000003b4
    );
  blk00000003_blk0000026d : XORCY
    port map (
      CI => blk00000003_sig000003af,
      LI => blk00000003_sig000003b0,
      O => blk00000003_sig000003b1
    );
  blk00000003_blk0000026c : XORCY
    port map (
      CI => blk00000003_sig000003ac,
      LI => blk00000003_sig000003ad,
      O => blk00000003_sig000003ae
    );
  blk00000003_blk0000026b : XORCY
    port map (
      CI => blk00000003_sig000003a9,
      LI => blk00000003_sig000003aa,
      O => blk00000003_sig000003ab
    );
  blk00000003_blk0000026a : XORCY
    port map (
      CI => blk00000003_sig000003a6,
      LI => blk00000003_sig000003a7,
      O => blk00000003_sig000003a8
    );
  blk00000003_blk00000269 : XORCY
    port map (
      CI => blk00000003_sig000003a3,
      LI => blk00000003_sig000003a4,
      O => blk00000003_sig000003a5
    );
  blk00000003_blk00000268 : XORCY
    port map (
      CI => blk00000003_sig000003a0,
      LI => blk00000003_sig000003a1,
      O => blk00000003_sig000003a2
    );
  blk00000003_blk00000267 : XORCY
    port map (
      CI => blk00000003_sig0000039d,
      LI => blk00000003_sig0000039e,
      O => blk00000003_sig0000039f
    );
  blk00000003_blk00000266 : XORCY
    port map (
      CI => blk00000003_sig0000039a,
      LI => blk00000003_sig0000039b,
      O => blk00000003_sig0000039c
    );
  blk00000003_blk00000265 : XORCY
    port map (
      CI => blk00000003_sig00000397,
      LI => blk00000003_sig00000398,
      O => blk00000003_sig00000399
    );
  blk00000003_blk00000264 : XORCY
    port map (
      CI => blk00000003_sig00000394,
      LI => blk00000003_sig00000395,
      O => blk00000003_sig00000396
    );
  blk00000003_blk00000263 : XORCY
    port map (
      CI => blk00000003_sig00000391,
      LI => blk00000003_sig00000392,
      O => blk00000003_sig00000393
    );
  blk00000003_blk00000262 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000038b,
      Q => blk00000003_sig00000390
    );
  blk00000003_blk00000261 : MUXCY
    port map (
      CI => blk00000003_sig0000038c,
      DI => blk00000003_sig0000038f,
      S => blk00000003_sig0000038d,
      O => blk00000003_sig00000378
    );
  blk00000003_blk00000260 : XORCY
    port map (
      CI => blk00000003_sig0000038c,
      LI => blk00000003_sig0000038d,
      O => blk00000003_sig0000038e
    );
  blk00000003_blk0000025f : MUXCY
    port map (
      CI => blk00000003_sig0000034b,
      DI => blk00000003_sig0000038a,
      S => blk00000003_sig0000034c,
      O => blk00000003_sig0000038b
    );
  blk00000003_blk0000025e : MUXCY
    port map (
      CI => blk00000003_sig00000378,
      DI => blk00000003_sig00000389,
      S => blk00000003_sig00000379,
      O => blk00000003_sig00000375
    );
  blk00000003_blk0000025d : MUXCY
    port map (
      CI => blk00000003_sig00000375,
      DI => blk00000003_sig00000388,
      S => blk00000003_sig00000376,
      O => blk00000003_sig00000372
    );
  blk00000003_blk0000025c : MUXCY
    port map (
      CI => blk00000003_sig00000372,
      DI => blk00000003_sig00000387,
      S => blk00000003_sig00000373,
      O => blk00000003_sig0000036f
    );
  blk00000003_blk0000025b : MUXCY
    port map (
      CI => blk00000003_sig0000036f,
      DI => blk00000003_sig00000386,
      S => blk00000003_sig00000370,
      O => blk00000003_sig0000036c
    );
  blk00000003_blk0000025a : MUXCY
    port map (
      CI => blk00000003_sig0000036c,
      DI => blk00000003_sig00000385,
      S => blk00000003_sig0000036d,
      O => blk00000003_sig00000369
    );
  blk00000003_blk00000259 : MUXCY
    port map (
      CI => blk00000003_sig00000369,
      DI => blk00000003_sig00000384,
      S => blk00000003_sig0000036a,
      O => blk00000003_sig00000366
    );
  blk00000003_blk00000258 : MUXCY
    port map (
      CI => blk00000003_sig00000366,
      DI => blk00000003_sig00000383,
      S => blk00000003_sig00000367,
      O => blk00000003_sig00000363
    );
  blk00000003_blk00000257 : MUXCY
    port map (
      CI => blk00000003_sig00000363,
      DI => blk00000003_sig00000382,
      S => blk00000003_sig00000364,
      O => blk00000003_sig00000360
    );
  blk00000003_blk00000256 : MUXCY
    port map (
      CI => blk00000003_sig00000360,
      DI => blk00000003_sig00000381,
      S => blk00000003_sig00000361,
      O => blk00000003_sig0000035d
    );
  blk00000003_blk00000255 : MUXCY
    port map (
      CI => blk00000003_sig0000035d,
      DI => blk00000003_sig00000380,
      S => blk00000003_sig0000035e,
      O => blk00000003_sig0000035a
    );
  blk00000003_blk00000254 : MUXCY
    port map (
      CI => blk00000003_sig0000035a,
      DI => blk00000003_sig0000037f,
      S => blk00000003_sig0000035b,
      O => blk00000003_sig00000357
    );
  blk00000003_blk00000253 : MUXCY
    port map (
      CI => blk00000003_sig00000357,
      DI => blk00000003_sig0000037e,
      S => blk00000003_sig00000358,
      O => blk00000003_sig00000354
    );
  blk00000003_blk00000252 : MUXCY
    port map (
      CI => blk00000003_sig00000354,
      DI => blk00000003_sig0000037d,
      S => blk00000003_sig00000355,
      O => blk00000003_sig00000351
    );
  blk00000003_blk00000251 : MUXCY
    port map (
      CI => blk00000003_sig00000351,
      DI => blk00000003_sig0000037c,
      S => blk00000003_sig00000352,
      O => blk00000003_sig0000034e
    );
  blk00000003_blk00000250 : MUXCY
    port map (
      CI => blk00000003_sig0000034e,
      DI => blk00000003_sig0000037b,
      S => blk00000003_sig0000034f,
      O => blk00000003_sig0000034b
    );
  blk00000003_blk0000024f : XORCY
    port map (
      CI => blk00000003_sig00000378,
      LI => blk00000003_sig00000379,
      O => blk00000003_sig0000037a
    );
  blk00000003_blk0000024e : XORCY
    port map (
      CI => blk00000003_sig00000375,
      LI => blk00000003_sig00000376,
      O => blk00000003_sig00000377
    );
  blk00000003_blk0000024d : XORCY
    port map (
      CI => blk00000003_sig00000372,
      LI => blk00000003_sig00000373,
      O => blk00000003_sig00000374
    );
  blk00000003_blk0000024c : XORCY
    port map (
      CI => blk00000003_sig0000036f,
      LI => blk00000003_sig00000370,
      O => blk00000003_sig00000371
    );
  blk00000003_blk0000024b : XORCY
    port map (
      CI => blk00000003_sig0000036c,
      LI => blk00000003_sig0000036d,
      O => blk00000003_sig0000036e
    );
  blk00000003_blk0000024a : XORCY
    port map (
      CI => blk00000003_sig00000369,
      LI => blk00000003_sig0000036a,
      O => blk00000003_sig0000036b
    );
  blk00000003_blk00000249 : XORCY
    port map (
      CI => blk00000003_sig00000366,
      LI => blk00000003_sig00000367,
      O => blk00000003_sig00000368
    );
  blk00000003_blk00000248 : XORCY
    port map (
      CI => blk00000003_sig00000363,
      LI => blk00000003_sig00000364,
      O => blk00000003_sig00000365
    );
  blk00000003_blk00000247 : XORCY
    port map (
      CI => blk00000003_sig00000360,
      LI => blk00000003_sig00000361,
      O => blk00000003_sig00000362
    );
  blk00000003_blk00000246 : XORCY
    port map (
      CI => blk00000003_sig0000035d,
      LI => blk00000003_sig0000035e,
      O => blk00000003_sig0000035f
    );
  blk00000003_blk00000245 : XORCY
    port map (
      CI => blk00000003_sig0000035a,
      LI => blk00000003_sig0000035b,
      O => blk00000003_sig0000035c
    );
  blk00000003_blk00000244 : XORCY
    port map (
      CI => blk00000003_sig00000357,
      LI => blk00000003_sig00000358,
      O => blk00000003_sig00000359
    );
  blk00000003_blk00000243 : XORCY
    port map (
      CI => blk00000003_sig00000354,
      LI => blk00000003_sig00000355,
      O => blk00000003_sig00000356
    );
  blk00000003_blk00000242 : XORCY
    port map (
      CI => blk00000003_sig00000351,
      LI => blk00000003_sig00000352,
      O => blk00000003_sig00000353
    );
  blk00000003_blk00000241 : XORCY
    port map (
      CI => blk00000003_sig0000034e,
      LI => blk00000003_sig0000034f,
      O => blk00000003_sig00000350
    );
  blk00000003_blk00000240 : XORCY
    port map (
      CI => blk00000003_sig0000034b,
      LI => blk00000003_sig0000034c,
      O => blk00000003_sig0000034d
    );
  blk00000003_blk0000023f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000345,
      Q => blk00000003_sig0000034a
    );
  blk00000003_blk0000023e : MUXCY
    port map (
      CI => blk00000003_sig00000346,
      DI => blk00000003_sig00000349,
      S => blk00000003_sig00000347,
      O => blk00000003_sig00000332
    );
  blk00000003_blk0000023d : XORCY
    port map (
      CI => blk00000003_sig00000346,
      LI => blk00000003_sig00000347,
      O => blk00000003_sig00000348
    );
  blk00000003_blk0000023c : MUXCY
    port map (
      CI => blk00000003_sig00000305,
      DI => blk00000003_sig00000344,
      S => blk00000003_sig00000306,
      O => blk00000003_sig00000345
    );
  blk00000003_blk0000023b : MUXCY
    port map (
      CI => blk00000003_sig00000332,
      DI => blk00000003_sig00000343,
      S => blk00000003_sig00000333,
      O => blk00000003_sig0000032f
    );
  blk00000003_blk0000023a : MUXCY
    port map (
      CI => blk00000003_sig0000032f,
      DI => blk00000003_sig00000342,
      S => blk00000003_sig00000330,
      O => blk00000003_sig0000032c
    );
  blk00000003_blk00000239 : MUXCY
    port map (
      CI => blk00000003_sig0000032c,
      DI => blk00000003_sig00000341,
      S => blk00000003_sig0000032d,
      O => blk00000003_sig00000329
    );
  blk00000003_blk00000238 : MUXCY
    port map (
      CI => blk00000003_sig00000329,
      DI => blk00000003_sig00000340,
      S => blk00000003_sig0000032a,
      O => blk00000003_sig00000326
    );
  blk00000003_blk00000237 : MUXCY
    port map (
      CI => blk00000003_sig00000326,
      DI => blk00000003_sig0000033f,
      S => blk00000003_sig00000327,
      O => blk00000003_sig00000323
    );
  blk00000003_blk00000236 : MUXCY
    port map (
      CI => blk00000003_sig00000323,
      DI => blk00000003_sig0000033e,
      S => blk00000003_sig00000324,
      O => blk00000003_sig00000320
    );
  blk00000003_blk00000235 : MUXCY
    port map (
      CI => blk00000003_sig00000320,
      DI => blk00000003_sig0000033d,
      S => blk00000003_sig00000321,
      O => blk00000003_sig0000031d
    );
  blk00000003_blk00000234 : MUXCY
    port map (
      CI => blk00000003_sig0000031d,
      DI => blk00000003_sig0000033c,
      S => blk00000003_sig0000031e,
      O => blk00000003_sig0000031a
    );
  blk00000003_blk00000233 : MUXCY
    port map (
      CI => blk00000003_sig0000031a,
      DI => blk00000003_sig0000033b,
      S => blk00000003_sig0000031b,
      O => blk00000003_sig00000317
    );
  blk00000003_blk00000232 : MUXCY
    port map (
      CI => blk00000003_sig00000317,
      DI => blk00000003_sig0000033a,
      S => blk00000003_sig00000318,
      O => blk00000003_sig00000314
    );
  blk00000003_blk00000231 : MUXCY
    port map (
      CI => blk00000003_sig00000314,
      DI => blk00000003_sig00000339,
      S => blk00000003_sig00000315,
      O => blk00000003_sig00000311
    );
  blk00000003_blk00000230 : MUXCY
    port map (
      CI => blk00000003_sig00000311,
      DI => blk00000003_sig00000338,
      S => blk00000003_sig00000312,
      O => blk00000003_sig0000030e
    );
  blk00000003_blk0000022f : MUXCY
    port map (
      CI => blk00000003_sig0000030e,
      DI => blk00000003_sig00000337,
      S => blk00000003_sig0000030f,
      O => blk00000003_sig0000030b
    );
  blk00000003_blk0000022e : MUXCY
    port map (
      CI => blk00000003_sig0000030b,
      DI => blk00000003_sig00000336,
      S => blk00000003_sig0000030c,
      O => blk00000003_sig00000308
    );
  blk00000003_blk0000022d : MUXCY
    port map (
      CI => blk00000003_sig00000308,
      DI => blk00000003_sig00000335,
      S => blk00000003_sig00000309,
      O => blk00000003_sig00000305
    );
  blk00000003_blk0000022c : XORCY
    port map (
      CI => blk00000003_sig00000332,
      LI => blk00000003_sig00000333,
      O => blk00000003_sig00000334
    );
  blk00000003_blk0000022b : XORCY
    port map (
      CI => blk00000003_sig0000032f,
      LI => blk00000003_sig00000330,
      O => blk00000003_sig00000331
    );
  blk00000003_blk0000022a : XORCY
    port map (
      CI => blk00000003_sig0000032c,
      LI => blk00000003_sig0000032d,
      O => blk00000003_sig0000032e
    );
  blk00000003_blk00000229 : XORCY
    port map (
      CI => blk00000003_sig00000329,
      LI => blk00000003_sig0000032a,
      O => blk00000003_sig0000032b
    );
  blk00000003_blk00000228 : XORCY
    port map (
      CI => blk00000003_sig00000326,
      LI => blk00000003_sig00000327,
      O => blk00000003_sig00000328
    );
  blk00000003_blk00000227 : XORCY
    port map (
      CI => blk00000003_sig00000323,
      LI => blk00000003_sig00000324,
      O => blk00000003_sig00000325
    );
  blk00000003_blk00000226 : XORCY
    port map (
      CI => blk00000003_sig00000320,
      LI => blk00000003_sig00000321,
      O => blk00000003_sig00000322
    );
  blk00000003_blk00000225 : XORCY
    port map (
      CI => blk00000003_sig0000031d,
      LI => blk00000003_sig0000031e,
      O => blk00000003_sig0000031f
    );
  blk00000003_blk00000224 : XORCY
    port map (
      CI => blk00000003_sig0000031a,
      LI => blk00000003_sig0000031b,
      O => blk00000003_sig0000031c
    );
  blk00000003_blk00000223 : XORCY
    port map (
      CI => blk00000003_sig00000317,
      LI => blk00000003_sig00000318,
      O => blk00000003_sig00000319
    );
  blk00000003_blk00000222 : XORCY
    port map (
      CI => blk00000003_sig00000314,
      LI => blk00000003_sig00000315,
      O => blk00000003_sig00000316
    );
  blk00000003_blk00000221 : XORCY
    port map (
      CI => blk00000003_sig00000311,
      LI => blk00000003_sig00000312,
      O => blk00000003_sig00000313
    );
  blk00000003_blk00000220 : XORCY
    port map (
      CI => blk00000003_sig0000030e,
      LI => blk00000003_sig0000030f,
      O => blk00000003_sig00000310
    );
  blk00000003_blk0000021f : XORCY
    port map (
      CI => blk00000003_sig0000030b,
      LI => blk00000003_sig0000030c,
      O => blk00000003_sig0000030d
    );
  blk00000003_blk0000021e : XORCY
    port map (
      CI => blk00000003_sig00000308,
      LI => blk00000003_sig00000309,
      O => blk00000003_sig0000030a
    );
  blk00000003_blk0000021d : XORCY
    port map (
      CI => blk00000003_sig00000305,
      LI => blk00000003_sig00000306,
      O => blk00000003_sig00000307
    );
  blk00000003_blk0000021c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002ff,
      Q => blk00000003_sig00000304
    );
  blk00000003_blk0000021b : MUXCY
    port map (
      CI => blk00000003_sig00000300,
      DI => blk00000003_sig00000303,
      S => blk00000003_sig00000301,
      O => blk00000003_sig000002ec
    );
  blk00000003_blk0000021a : XORCY
    port map (
      CI => blk00000003_sig00000300,
      LI => blk00000003_sig00000301,
      O => blk00000003_sig00000302
    );
  blk00000003_blk00000219 : MUXCY
    port map (
      CI => blk00000003_sig000002bf,
      DI => blk00000003_sig000002fe,
      S => blk00000003_sig000002c0,
      O => blk00000003_sig000002ff
    );
  blk00000003_blk00000218 : MUXCY
    port map (
      CI => blk00000003_sig000002ec,
      DI => blk00000003_sig000002fd,
      S => blk00000003_sig000002ed,
      O => blk00000003_sig000002e9
    );
  blk00000003_blk00000217 : MUXCY
    port map (
      CI => blk00000003_sig000002e9,
      DI => blk00000003_sig000002fc,
      S => blk00000003_sig000002ea,
      O => blk00000003_sig000002e6
    );
  blk00000003_blk00000216 : MUXCY
    port map (
      CI => blk00000003_sig000002e6,
      DI => blk00000003_sig000002fb,
      S => blk00000003_sig000002e7,
      O => blk00000003_sig000002e3
    );
  blk00000003_blk00000215 : MUXCY
    port map (
      CI => blk00000003_sig000002e3,
      DI => blk00000003_sig000002fa,
      S => blk00000003_sig000002e4,
      O => blk00000003_sig000002e0
    );
  blk00000003_blk00000214 : MUXCY
    port map (
      CI => blk00000003_sig000002e0,
      DI => blk00000003_sig000002f9,
      S => blk00000003_sig000002e1,
      O => blk00000003_sig000002dd
    );
  blk00000003_blk00000213 : MUXCY
    port map (
      CI => blk00000003_sig000002dd,
      DI => blk00000003_sig000002f8,
      S => blk00000003_sig000002de,
      O => blk00000003_sig000002da
    );
  blk00000003_blk00000212 : MUXCY
    port map (
      CI => blk00000003_sig000002da,
      DI => blk00000003_sig000002f7,
      S => blk00000003_sig000002db,
      O => blk00000003_sig000002d7
    );
  blk00000003_blk00000211 : MUXCY
    port map (
      CI => blk00000003_sig000002d7,
      DI => blk00000003_sig000002f6,
      S => blk00000003_sig000002d8,
      O => blk00000003_sig000002d4
    );
  blk00000003_blk00000210 : MUXCY
    port map (
      CI => blk00000003_sig000002d4,
      DI => blk00000003_sig000002f5,
      S => blk00000003_sig000002d5,
      O => blk00000003_sig000002d1
    );
  blk00000003_blk0000020f : MUXCY
    port map (
      CI => blk00000003_sig000002d1,
      DI => blk00000003_sig000002f4,
      S => blk00000003_sig000002d2,
      O => blk00000003_sig000002ce
    );
  blk00000003_blk0000020e : MUXCY
    port map (
      CI => blk00000003_sig000002ce,
      DI => blk00000003_sig000002f3,
      S => blk00000003_sig000002cf,
      O => blk00000003_sig000002cb
    );
  blk00000003_blk0000020d : MUXCY
    port map (
      CI => blk00000003_sig000002cb,
      DI => blk00000003_sig000002f2,
      S => blk00000003_sig000002cc,
      O => blk00000003_sig000002c8
    );
  blk00000003_blk0000020c : MUXCY
    port map (
      CI => blk00000003_sig000002c8,
      DI => blk00000003_sig000002f1,
      S => blk00000003_sig000002c9,
      O => blk00000003_sig000002c5
    );
  blk00000003_blk0000020b : MUXCY
    port map (
      CI => blk00000003_sig000002c5,
      DI => blk00000003_sig000002f0,
      S => blk00000003_sig000002c6,
      O => blk00000003_sig000002c2
    );
  blk00000003_blk0000020a : MUXCY
    port map (
      CI => blk00000003_sig000002c2,
      DI => blk00000003_sig000002ef,
      S => blk00000003_sig000002c3,
      O => blk00000003_sig000002bf
    );
  blk00000003_blk00000209 : XORCY
    port map (
      CI => blk00000003_sig000002ec,
      LI => blk00000003_sig000002ed,
      O => blk00000003_sig000002ee
    );
  blk00000003_blk00000208 : XORCY
    port map (
      CI => blk00000003_sig000002e9,
      LI => blk00000003_sig000002ea,
      O => blk00000003_sig000002eb
    );
  blk00000003_blk00000207 : XORCY
    port map (
      CI => blk00000003_sig000002e6,
      LI => blk00000003_sig000002e7,
      O => blk00000003_sig000002e8
    );
  blk00000003_blk00000206 : XORCY
    port map (
      CI => blk00000003_sig000002e3,
      LI => blk00000003_sig000002e4,
      O => blk00000003_sig000002e5
    );
  blk00000003_blk00000205 : XORCY
    port map (
      CI => blk00000003_sig000002e0,
      LI => blk00000003_sig000002e1,
      O => blk00000003_sig000002e2
    );
  blk00000003_blk00000204 : XORCY
    port map (
      CI => blk00000003_sig000002dd,
      LI => blk00000003_sig000002de,
      O => blk00000003_sig000002df
    );
  blk00000003_blk00000203 : XORCY
    port map (
      CI => blk00000003_sig000002da,
      LI => blk00000003_sig000002db,
      O => blk00000003_sig000002dc
    );
  blk00000003_blk00000202 : XORCY
    port map (
      CI => blk00000003_sig000002d7,
      LI => blk00000003_sig000002d8,
      O => blk00000003_sig000002d9
    );
  blk00000003_blk00000201 : XORCY
    port map (
      CI => blk00000003_sig000002d4,
      LI => blk00000003_sig000002d5,
      O => blk00000003_sig000002d6
    );
  blk00000003_blk00000200 : XORCY
    port map (
      CI => blk00000003_sig000002d1,
      LI => blk00000003_sig000002d2,
      O => blk00000003_sig000002d3
    );
  blk00000003_blk000001ff : XORCY
    port map (
      CI => blk00000003_sig000002ce,
      LI => blk00000003_sig000002cf,
      O => blk00000003_sig000002d0
    );
  blk00000003_blk000001fe : XORCY
    port map (
      CI => blk00000003_sig000002cb,
      LI => blk00000003_sig000002cc,
      O => blk00000003_sig000002cd
    );
  blk00000003_blk000001fd : XORCY
    port map (
      CI => blk00000003_sig000002c8,
      LI => blk00000003_sig000002c9,
      O => blk00000003_sig000002ca
    );
  blk00000003_blk000001fc : XORCY
    port map (
      CI => blk00000003_sig000002c5,
      LI => blk00000003_sig000002c6,
      O => blk00000003_sig000002c7
    );
  blk00000003_blk000001fb : XORCY
    port map (
      CI => blk00000003_sig000002c2,
      LI => blk00000003_sig000002c3,
      O => blk00000003_sig000002c4
    );
  blk00000003_blk000001fa : XORCY
    port map (
      CI => blk00000003_sig000002bf,
      LI => blk00000003_sig000002c0,
      O => blk00000003_sig000002c1
    );
  blk00000003_blk000001f9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002b9,
      Q => blk00000003_sig000002be
    );
  blk00000003_blk000001f8 : MUXCY
    port map (
      CI => blk00000003_sig000002ba,
      DI => blk00000003_sig000002bd,
      S => blk00000003_sig000002bb,
      O => blk00000003_sig000002a6
    );
  blk00000003_blk000001f7 : XORCY
    port map (
      CI => blk00000003_sig000002ba,
      LI => blk00000003_sig000002bb,
      O => blk00000003_sig000002bc
    );
  blk00000003_blk000001f6 : MUXCY
    port map (
      CI => blk00000003_sig00000279,
      DI => blk00000003_sig000002b8,
      S => blk00000003_sig0000027a,
      O => blk00000003_sig000002b9
    );
  blk00000003_blk000001f5 : MUXCY
    port map (
      CI => blk00000003_sig000002a6,
      DI => blk00000003_sig000002b7,
      S => blk00000003_sig000002a7,
      O => blk00000003_sig000002a3
    );
  blk00000003_blk000001f4 : MUXCY
    port map (
      CI => blk00000003_sig000002a3,
      DI => blk00000003_sig000002b6,
      S => blk00000003_sig000002a4,
      O => blk00000003_sig000002a0
    );
  blk00000003_blk000001f3 : MUXCY
    port map (
      CI => blk00000003_sig000002a0,
      DI => blk00000003_sig000002b5,
      S => blk00000003_sig000002a1,
      O => blk00000003_sig0000029d
    );
  blk00000003_blk000001f2 : MUXCY
    port map (
      CI => blk00000003_sig0000029d,
      DI => blk00000003_sig000002b4,
      S => blk00000003_sig0000029e,
      O => blk00000003_sig0000029a
    );
  blk00000003_blk000001f1 : MUXCY
    port map (
      CI => blk00000003_sig0000029a,
      DI => blk00000003_sig000002b3,
      S => blk00000003_sig0000029b,
      O => blk00000003_sig00000297
    );
  blk00000003_blk000001f0 : MUXCY
    port map (
      CI => blk00000003_sig00000297,
      DI => blk00000003_sig000002b2,
      S => blk00000003_sig00000298,
      O => blk00000003_sig00000294
    );
  blk00000003_blk000001ef : MUXCY
    port map (
      CI => blk00000003_sig00000294,
      DI => blk00000003_sig000002b1,
      S => blk00000003_sig00000295,
      O => blk00000003_sig00000291
    );
  blk00000003_blk000001ee : MUXCY
    port map (
      CI => blk00000003_sig00000291,
      DI => blk00000003_sig000002b0,
      S => blk00000003_sig00000292,
      O => blk00000003_sig0000028e
    );
  blk00000003_blk000001ed : MUXCY
    port map (
      CI => blk00000003_sig0000028e,
      DI => blk00000003_sig000002af,
      S => blk00000003_sig0000028f,
      O => blk00000003_sig0000028b
    );
  blk00000003_blk000001ec : MUXCY
    port map (
      CI => blk00000003_sig0000028b,
      DI => blk00000003_sig000002ae,
      S => blk00000003_sig0000028c,
      O => blk00000003_sig00000288
    );
  blk00000003_blk000001eb : MUXCY
    port map (
      CI => blk00000003_sig00000288,
      DI => blk00000003_sig000002ad,
      S => blk00000003_sig00000289,
      O => blk00000003_sig00000285
    );
  blk00000003_blk000001ea : MUXCY
    port map (
      CI => blk00000003_sig00000285,
      DI => blk00000003_sig000002ac,
      S => blk00000003_sig00000286,
      O => blk00000003_sig00000282
    );
  blk00000003_blk000001e9 : MUXCY
    port map (
      CI => blk00000003_sig00000282,
      DI => blk00000003_sig000002ab,
      S => blk00000003_sig00000283,
      O => blk00000003_sig0000027f
    );
  blk00000003_blk000001e8 : MUXCY
    port map (
      CI => blk00000003_sig0000027f,
      DI => blk00000003_sig000002aa,
      S => blk00000003_sig00000280,
      O => blk00000003_sig0000027c
    );
  blk00000003_blk000001e7 : MUXCY
    port map (
      CI => blk00000003_sig0000027c,
      DI => blk00000003_sig000002a9,
      S => blk00000003_sig0000027d,
      O => blk00000003_sig00000279
    );
  blk00000003_blk000001e6 : XORCY
    port map (
      CI => blk00000003_sig000002a6,
      LI => blk00000003_sig000002a7,
      O => blk00000003_sig000002a8
    );
  blk00000003_blk000001e5 : XORCY
    port map (
      CI => blk00000003_sig000002a3,
      LI => blk00000003_sig000002a4,
      O => blk00000003_sig000002a5
    );
  blk00000003_blk000001e4 : XORCY
    port map (
      CI => blk00000003_sig000002a0,
      LI => blk00000003_sig000002a1,
      O => blk00000003_sig000002a2
    );
  blk00000003_blk000001e3 : XORCY
    port map (
      CI => blk00000003_sig0000029d,
      LI => blk00000003_sig0000029e,
      O => blk00000003_sig0000029f
    );
  blk00000003_blk000001e2 : XORCY
    port map (
      CI => blk00000003_sig0000029a,
      LI => blk00000003_sig0000029b,
      O => blk00000003_sig0000029c
    );
  blk00000003_blk000001e1 : XORCY
    port map (
      CI => blk00000003_sig00000297,
      LI => blk00000003_sig00000298,
      O => blk00000003_sig00000299
    );
  blk00000003_blk000001e0 : XORCY
    port map (
      CI => blk00000003_sig00000294,
      LI => blk00000003_sig00000295,
      O => blk00000003_sig00000296
    );
  blk00000003_blk000001df : XORCY
    port map (
      CI => blk00000003_sig00000291,
      LI => blk00000003_sig00000292,
      O => blk00000003_sig00000293
    );
  blk00000003_blk000001de : XORCY
    port map (
      CI => blk00000003_sig0000028e,
      LI => blk00000003_sig0000028f,
      O => blk00000003_sig00000290
    );
  blk00000003_blk000001dd : XORCY
    port map (
      CI => blk00000003_sig0000028b,
      LI => blk00000003_sig0000028c,
      O => blk00000003_sig0000028d
    );
  blk00000003_blk000001dc : XORCY
    port map (
      CI => blk00000003_sig00000288,
      LI => blk00000003_sig00000289,
      O => blk00000003_sig0000028a
    );
  blk00000003_blk000001db : XORCY
    port map (
      CI => blk00000003_sig00000285,
      LI => blk00000003_sig00000286,
      O => blk00000003_sig00000287
    );
  blk00000003_blk000001da : XORCY
    port map (
      CI => blk00000003_sig00000282,
      LI => blk00000003_sig00000283,
      O => blk00000003_sig00000284
    );
  blk00000003_blk000001d9 : XORCY
    port map (
      CI => blk00000003_sig0000027f,
      LI => blk00000003_sig00000280,
      O => blk00000003_sig00000281
    );
  blk00000003_blk000001d8 : XORCY
    port map (
      CI => blk00000003_sig0000027c,
      LI => blk00000003_sig0000027d,
      O => blk00000003_sig0000027e
    );
  blk00000003_blk000001d7 : XORCY
    port map (
      CI => blk00000003_sig00000279,
      LI => blk00000003_sig0000027a,
      O => blk00000003_sig0000027b
    );
  blk00000003_blk000001d6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000273,
      Q => blk00000003_sig00000278
    );
  blk00000003_blk000001d5 : MUXCY
    port map (
      CI => blk00000003_sig00000274,
      DI => blk00000003_sig00000277,
      S => blk00000003_sig00000275,
      O => blk00000003_sig00000260
    );
  blk00000003_blk000001d4 : XORCY
    port map (
      CI => blk00000003_sig00000274,
      LI => blk00000003_sig00000275,
      O => blk00000003_sig00000276
    );
  blk00000003_blk000001d3 : MUXCY
    port map (
      CI => blk00000003_sig00000233,
      DI => blk00000003_sig00000272,
      S => blk00000003_sig00000234,
      O => blk00000003_sig00000273
    );
  blk00000003_blk000001d2 : MUXCY
    port map (
      CI => blk00000003_sig00000260,
      DI => blk00000003_sig00000271,
      S => blk00000003_sig00000261,
      O => blk00000003_sig0000025d
    );
  blk00000003_blk000001d1 : MUXCY
    port map (
      CI => blk00000003_sig0000025d,
      DI => blk00000003_sig00000270,
      S => blk00000003_sig0000025e,
      O => blk00000003_sig0000025a
    );
  blk00000003_blk000001d0 : MUXCY
    port map (
      CI => blk00000003_sig0000025a,
      DI => blk00000003_sig0000026f,
      S => blk00000003_sig0000025b,
      O => blk00000003_sig00000257
    );
  blk00000003_blk000001cf : MUXCY
    port map (
      CI => blk00000003_sig00000257,
      DI => blk00000003_sig0000026e,
      S => blk00000003_sig00000258,
      O => blk00000003_sig00000254
    );
  blk00000003_blk000001ce : MUXCY
    port map (
      CI => blk00000003_sig00000254,
      DI => blk00000003_sig0000026d,
      S => blk00000003_sig00000255,
      O => blk00000003_sig00000251
    );
  blk00000003_blk000001cd : MUXCY
    port map (
      CI => blk00000003_sig00000251,
      DI => blk00000003_sig0000026c,
      S => blk00000003_sig00000252,
      O => blk00000003_sig0000024e
    );
  blk00000003_blk000001cc : MUXCY
    port map (
      CI => blk00000003_sig0000024e,
      DI => blk00000003_sig0000026b,
      S => blk00000003_sig0000024f,
      O => blk00000003_sig0000024b
    );
  blk00000003_blk000001cb : MUXCY
    port map (
      CI => blk00000003_sig0000024b,
      DI => blk00000003_sig0000026a,
      S => blk00000003_sig0000024c,
      O => blk00000003_sig00000248
    );
  blk00000003_blk000001ca : MUXCY
    port map (
      CI => blk00000003_sig00000248,
      DI => blk00000003_sig00000269,
      S => blk00000003_sig00000249,
      O => blk00000003_sig00000245
    );
  blk00000003_blk000001c9 : MUXCY
    port map (
      CI => blk00000003_sig00000245,
      DI => blk00000003_sig00000268,
      S => blk00000003_sig00000246,
      O => blk00000003_sig00000242
    );
  blk00000003_blk000001c8 : MUXCY
    port map (
      CI => blk00000003_sig00000242,
      DI => blk00000003_sig00000267,
      S => blk00000003_sig00000243,
      O => blk00000003_sig0000023f
    );
  blk00000003_blk000001c7 : MUXCY
    port map (
      CI => blk00000003_sig0000023f,
      DI => blk00000003_sig00000266,
      S => blk00000003_sig00000240,
      O => blk00000003_sig0000023c
    );
  blk00000003_blk000001c6 : MUXCY
    port map (
      CI => blk00000003_sig0000023c,
      DI => blk00000003_sig00000265,
      S => blk00000003_sig0000023d,
      O => blk00000003_sig00000239
    );
  blk00000003_blk000001c5 : MUXCY
    port map (
      CI => blk00000003_sig00000239,
      DI => blk00000003_sig00000264,
      S => blk00000003_sig0000023a,
      O => blk00000003_sig00000236
    );
  blk00000003_blk000001c4 : MUXCY
    port map (
      CI => blk00000003_sig00000236,
      DI => blk00000003_sig00000263,
      S => blk00000003_sig00000237,
      O => blk00000003_sig00000233
    );
  blk00000003_blk000001c3 : XORCY
    port map (
      CI => blk00000003_sig00000260,
      LI => blk00000003_sig00000261,
      O => blk00000003_sig00000262
    );
  blk00000003_blk000001c2 : XORCY
    port map (
      CI => blk00000003_sig0000025d,
      LI => blk00000003_sig0000025e,
      O => blk00000003_sig0000025f
    );
  blk00000003_blk000001c1 : XORCY
    port map (
      CI => blk00000003_sig0000025a,
      LI => blk00000003_sig0000025b,
      O => blk00000003_sig0000025c
    );
  blk00000003_blk000001c0 : XORCY
    port map (
      CI => blk00000003_sig00000257,
      LI => blk00000003_sig00000258,
      O => blk00000003_sig00000259
    );
  blk00000003_blk000001bf : XORCY
    port map (
      CI => blk00000003_sig00000254,
      LI => blk00000003_sig00000255,
      O => blk00000003_sig00000256
    );
  blk00000003_blk000001be : XORCY
    port map (
      CI => blk00000003_sig00000251,
      LI => blk00000003_sig00000252,
      O => blk00000003_sig00000253
    );
  blk00000003_blk000001bd : XORCY
    port map (
      CI => blk00000003_sig0000024e,
      LI => blk00000003_sig0000024f,
      O => blk00000003_sig00000250
    );
  blk00000003_blk000001bc : XORCY
    port map (
      CI => blk00000003_sig0000024b,
      LI => blk00000003_sig0000024c,
      O => blk00000003_sig0000024d
    );
  blk00000003_blk000001bb : XORCY
    port map (
      CI => blk00000003_sig00000248,
      LI => blk00000003_sig00000249,
      O => blk00000003_sig0000024a
    );
  blk00000003_blk000001ba : XORCY
    port map (
      CI => blk00000003_sig00000245,
      LI => blk00000003_sig00000246,
      O => blk00000003_sig00000247
    );
  blk00000003_blk000001b9 : XORCY
    port map (
      CI => blk00000003_sig00000242,
      LI => blk00000003_sig00000243,
      O => blk00000003_sig00000244
    );
  blk00000003_blk000001b8 : XORCY
    port map (
      CI => blk00000003_sig0000023f,
      LI => blk00000003_sig00000240,
      O => blk00000003_sig00000241
    );
  blk00000003_blk000001b7 : XORCY
    port map (
      CI => blk00000003_sig0000023c,
      LI => blk00000003_sig0000023d,
      O => blk00000003_sig0000023e
    );
  blk00000003_blk000001b6 : XORCY
    port map (
      CI => blk00000003_sig00000239,
      LI => blk00000003_sig0000023a,
      O => blk00000003_sig0000023b
    );
  blk00000003_blk000001b5 : XORCY
    port map (
      CI => blk00000003_sig00000236,
      LI => blk00000003_sig00000237,
      O => blk00000003_sig00000238
    );
  blk00000003_blk000001b4 : XORCY
    port map (
      CI => blk00000003_sig00000233,
      LI => blk00000003_sig00000234,
      O => blk00000003_sig00000235
    );
  blk00000003_blk000001b3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000022d,
      Q => blk00000003_sig00000232
    );
  blk00000003_blk000001b2 : MUXCY
    port map (
      CI => blk00000003_sig0000022e,
      DI => blk00000003_sig00000231,
      S => blk00000003_sig0000022f,
      O => blk00000003_sig0000021a
    );
  blk00000003_blk000001b1 : XORCY
    port map (
      CI => blk00000003_sig0000022e,
      LI => blk00000003_sig0000022f,
      O => blk00000003_sig00000230
    );
  blk00000003_blk000001b0 : MUXCY
    port map (
      CI => blk00000003_sig000001ed,
      DI => blk00000003_sig0000022c,
      S => blk00000003_sig000001ee,
      O => blk00000003_sig0000022d
    );
  blk00000003_blk000001af : MUXCY
    port map (
      CI => blk00000003_sig0000021a,
      DI => blk00000003_sig0000022b,
      S => blk00000003_sig0000021b,
      O => blk00000003_sig00000217
    );
  blk00000003_blk000001ae : MUXCY
    port map (
      CI => blk00000003_sig00000217,
      DI => blk00000003_sig0000022a,
      S => blk00000003_sig00000218,
      O => blk00000003_sig00000214
    );
  blk00000003_blk000001ad : MUXCY
    port map (
      CI => blk00000003_sig00000214,
      DI => blk00000003_sig00000229,
      S => blk00000003_sig00000215,
      O => blk00000003_sig00000211
    );
  blk00000003_blk000001ac : MUXCY
    port map (
      CI => blk00000003_sig00000211,
      DI => blk00000003_sig00000228,
      S => blk00000003_sig00000212,
      O => blk00000003_sig0000020e
    );
  blk00000003_blk000001ab : MUXCY
    port map (
      CI => blk00000003_sig0000020e,
      DI => blk00000003_sig00000227,
      S => blk00000003_sig0000020f,
      O => blk00000003_sig0000020b
    );
  blk00000003_blk000001aa : MUXCY
    port map (
      CI => blk00000003_sig0000020b,
      DI => blk00000003_sig00000226,
      S => blk00000003_sig0000020c,
      O => blk00000003_sig00000208
    );
  blk00000003_blk000001a9 : MUXCY
    port map (
      CI => blk00000003_sig00000208,
      DI => blk00000003_sig00000225,
      S => blk00000003_sig00000209,
      O => blk00000003_sig00000205
    );
  blk00000003_blk000001a8 : MUXCY
    port map (
      CI => blk00000003_sig00000205,
      DI => blk00000003_sig00000224,
      S => blk00000003_sig00000206,
      O => blk00000003_sig00000202
    );
  blk00000003_blk000001a7 : MUXCY
    port map (
      CI => blk00000003_sig00000202,
      DI => blk00000003_sig00000223,
      S => blk00000003_sig00000203,
      O => blk00000003_sig000001ff
    );
  blk00000003_blk000001a6 : MUXCY
    port map (
      CI => blk00000003_sig000001ff,
      DI => blk00000003_sig00000222,
      S => blk00000003_sig00000200,
      O => blk00000003_sig000001fc
    );
  blk00000003_blk000001a5 : MUXCY
    port map (
      CI => blk00000003_sig000001fc,
      DI => blk00000003_sig00000221,
      S => blk00000003_sig000001fd,
      O => blk00000003_sig000001f9
    );
  blk00000003_blk000001a4 : MUXCY
    port map (
      CI => blk00000003_sig000001f9,
      DI => blk00000003_sig00000220,
      S => blk00000003_sig000001fa,
      O => blk00000003_sig000001f6
    );
  blk00000003_blk000001a3 : MUXCY
    port map (
      CI => blk00000003_sig000001f6,
      DI => blk00000003_sig0000021f,
      S => blk00000003_sig000001f7,
      O => blk00000003_sig000001f3
    );
  blk00000003_blk000001a2 : MUXCY
    port map (
      CI => blk00000003_sig000001f3,
      DI => blk00000003_sig0000021e,
      S => blk00000003_sig000001f4,
      O => blk00000003_sig000001f0
    );
  blk00000003_blk000001a1 : MUXCY
    port map (
      CI => blk00000003_sig000001f0,
      DI => blk00000003_sig0000021d,
      S => blk00000003_sig000001f1,
      O => blk00000003_sig000001ed
    );
  blk00000003_blk000001a0 : XORCY
    port map (
      CI => blk00000003_sig0000021a,
      LI => blk00000003_sig0000021b,
      O => blk00000003_sig0000021c
    );
  blk00000003_blk0000019f : XORCY
    port map (
      CI => blk00000003_sig00000217,
      LI => blk00000003_sig00000218,
      O => blk00000003_sig00000219
    );
  blk00000003_blk0000019e : XORCY
    port map (
      CI => blk00000003_sig00000214,
      LI => blk00000003_sig00000215,
      O => blk00000003_sig00000216
    );
  blk00000003_blk0000019d : XORCY
    port map (
      CI => blk00000003_sig00000211,
      LI => blk00000003_sig00000212,
      O => blk00000003_sig00000213
    );
  blk00000003_blk0000019c : XORCY
    port map (
      CI => blk00000003_sig0000020e,
      LI => blk00000003_sig0000020f,
      O => blk00000003_sig00000210
    );
  blk00000003_blk0000019b : XORCY
    port map (
      CI => blk00000003_sig0000020b,
      LI => blk00000003_sig0000020c,
      O => blk00000003_sig0000020d
    );
  blk00000003_blk0000019a : XORCY
    port map (
      CI => blk00000003_sig00000208,
      LI => blk00000003_sig00000209,
      O => blk00000003_sig0000020a
    );
  blk00000003_blk00000199 : XORCY
    port map (
      CI => blk00000003_sig00000205,
      LI => blk00000003_sig00000206,
      O => blk00000003_sig00000207
    );
  blk00000003_blk00000198 : XORCY
    port map (
      CI => blk00000003_sig00000202,
      LI => blk00000003_sig00000203,
      O => blk00000003_sig00000204
    );
  blk00000003_blk00000197 : XORCY
    port map (
      CI => blk00000003_sig000001ff,
      LI => blk00000003_sig00000200,
      O => blk00000003_sig00000201
    );
  blk00000003_blk00000196 : XORCY
    port map (
      CI => blk00000003_sig000001fc,
      LI => blk00000003_sig000001fd,
      O => blk00000003_sig000001fe
    );
  blk00000003_blk00000195 : XORCY
    port map (
      CI => blk00000003_sig000001f9,
      LI => blk00000003_sig000001fa,
      O => blk00000003_sig000001fb
    );
  blk00000003_blk00000194 : XORCY
    port map (
      CI => blk00000003_sig000001f6,
      LI => blk00000003_sig000001f7,
      O => blk00000003_sig000001f8
    );
  blk00000003_blk00000193 : XORCY
    port map (
      CI => blk00000003_sig000001f3,
      LI => blk00000003_sig000001f4,
      O => blk00000003_sig000001f5
    );
  blk00000003_blk00000192 : XORCY
    port map (
      CI => blk00000003_sig000001f0,
      LI => blk00000003_sig000001f1,
      O => blk00000003_sig000001f2
    );
  blk00000003_blk00000191 : XORCY
    port map (
      CI => blk00000003_sig000001ed,
      LI => blk00000003_sig000001ee,
      O => blk00000003_sig000001ef
    );
  blk00000003_blk00000190 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001e9,
      Q => blk00000003_sig000001ec
    );
  blk00000003_blk0000018f : MUXCY
    port map (
      CI => NlwRenamedSig_OI_rfd,
      DI => blk00000003_sig0000009b,
      S => blk00000003_sig000001ea,
      O => blk00000003_sig000001e6
    );
  blk00000003_blk0000018e : XORCY
    port map (
      CI => NlwRenamedSig_OI_rfd,
      LI => blk00000003_sig000001ea,
      O => blk00000003_sig000001eb
    );
  blk00000003_blk0000018d : MUXCY
    port map (
      CI => blk00000003_sig000001bb,
      DI => blk00000003_sig00000043,
      S => NlwRenamedSig_OI_rfd,
      O => blk00000003_sig000001e9
    );
  blk00000003_blk0000018c : MUXCY
    port map (
      CI => blk00000003_sig000001e6,
      DI => blk00000003_sig00000043,
      S => blk00000003_sig000001e7,
      O => blk00000003_sig000001e3
    );
  blk00000003_blk0000018b : MUXCY
    port map (
      CI => blk00000003_sig000001e3,
      DI => blk00000003_sig00000043,
      S => blk00000003_sig000001e4,
      O => blk00000003_sig000001e0
    );
  blk00000003_blk0000018a : MUXCY
    port map (
      CI => blk00000003_sig000001e0,
      DI => blk00000003_sig00000043,
      S => blk00000003_sig000001e1,
      O => blk00000003_sig000001dd
    );
  blk00000003_blk00000189 : MUXCY
    port map (
      CI => blk00000003_sig000001dd,
      DI => blk00000003_sig00000043,
      S => blk00000003_sig000001de,
      O => blk00000003_sig000001da
    );
  blk00000003_blk00000188 : MUXCY
    port map (
      CI => blk00000003_sig000001da,
      DI => blk00000003_sig00000043,
      S => blk00000003_sig000001db,
      O => blk00000003_sig000001d7
    );
  blk00000003_blk00000187 : MUXCY
    port map (
      CI => blk00000003_sig000001d7,
      DI => blk00000003_sig00000043,
      S => blk00000003_sig000001d8,
      O => blk00000003_sig000001d4
    );
  blk00000003_blk00000186 : MUXCY
    port map (
      CI => blk00000003_sig000001d4,
      DI => blk00000003_sig00000043,
      S => blk00000003_sig000001d5,
      O => blk00000003_sig000001d1
    );
  blk00000003_blk00000185 : MUXCY
    port map (
      CI => blk00000003_sig000001d1,
      DI => blk00000003_sig00000043,
      S => blk00000003_sig000001d2,
      O => blk00000003_sig000001ce
    );
  blk00000003_blk00000184 : MUXCY
    port map (
      CI => blk00000003_sig000001ce,
      DI => blk00000003_sig00000043,
      S => blk00000003_sig000001cf,
      O => blk00000003_sig000001cb
    );
  blk00000003_blk00000183 : MUXCY
    port map (
      CI => blk00000003_sig000001cb,
      DI => blk00000003_sig00000043,
      S => blk00000003_sig000001cc,
      O => blk00000003_sig000001c8
    );
  blk00000003_blk00000182 : MUXCY
    port map (
      CI => blk00000003_sig000001c8,
      DI => blk00000003_sig00000043,
      S => blk00000003_sig000001c9,
      O => blk00000003_sig000001c5
    );
  blk00000003_blk00000181 : MUXCY
    port map (
      CI => blk00000003_sig000001c5,
      DI => blk00000003_sig00000043,
      S => blk00000003_sig000001c6,
      O => blk00000003_sig000001c2
    );
  blk00000003_blk00000180 : MUXCY
    port map (
      CI => blk00000003_sig000001c2,
      DI => blk00000003_sig00000043,
      S => blk00000003_sig000001c3,
      O => blk00000003_sig000001bf
    );
  blk00000003_blk0000017f : MUXCY
    port map (
      CI => blk00000003_sig000001bf,
      DI => blk00000003_sig00000043,
      S => blk00000003_sig000001c0,
      O => blk00000003_sig000001bc
    );
  blk00000003_blk0000017e : MUXCY
    port map (
      CI => blk00000003_sig000001bc,
      DI => blk00000003_sig00000043,
      S => blk00000003_sig000001bd,
      O => blk00000003_sig000001bb
    );
  blk00000003_blk0000017d : XORCY
    port map (
      CI => blk00000003_sig000001e6,
      LI => blk00000003_sig000001e7,
      O => blk00000003_sig000001e8
    );
  blk00000003_blk0000017c : XORCY
    port map (
      CI => blk00000003_sig000001e3,
      LI => blk00000003_sig000001e4,
      O => blk00000003_sig000001e5
    );
  blk00000003_blk0000017b : XORCY
    port map (
      CI => blk00000003_sig000001e0,
      LI => blk00000003_sig000001e1,
      O => blk00000003_sig000001e2
    );
  blk00000003_blk0000017a : XORCY
    port map (
      CI => blk00000003_sig000001dd,
      LI => blk00000003_sig000001de,
      O => blk00000003_sig000001df
    );
  blk00000003_blk00000179 : XORCY
    port map (
      CI => blk00000003_sig000001da,
      LI => blk00000003_sig000001db,
      O => blk00000003_sig000001dc
    );
  blk00000003_blk00000178 : XORCY
    port map (
      CI => blk00000003_sig000001d7,
      LI => blk00000003_sig000001d8,
      O => blk00000003_sig000001d9
    );
  blk00000003_blk00000177 : XORCY
    port map (
      CI => blk00000003_sig000001d4,
      LI => blk00000003_sig000001d5,
      O => blk00000003_sig000001d6
    );
  blk00000003_blk00000176 : XORCY
    port map (
      CI => blk00000003_sig000001d1,
      LI => blk00000003_sig000001d2,
      O => blk00000003_sig000001d3
    );
  blk00000003_blk00000175 : XORCY
    port map (
      CI => blk00000003_sig000001ce,
      LI => blk00000003_sig000001cf,
      O => blk00000003_sig000001d0
    );
  blk00000003_blk00000174 : XORCY
    port map (
      CI => blk00000003_sig000001cb,
      LI => blk00000003_sig000001cc,
      O => blk00000003_sig000001cd
    );
  blk00000003_blk00000173 : XORCY
    port map (
      CI => blk00000003_sig000001c8,
      LI => blk00000003_sig000001c9,
      O => blk00000003_sig000001ca
    );
  blk00000003_blk00000172 : XORCY
    port map (
      CI => blk00000003_sig000001c5,
      LI => blk00000003_sig000001c6,
      O => blk00000003_sig000001c7
    );
  blk00000003_blk00000171 : XORCY
    port map (
      CI => blk00000003_sig000001c2,
      LI => blk00000003_sig000001c3,
      O => blk00000003_sig000001c4
    );
  blk00000003_blk00000170 : XORCY
    port map (
      CI => blk00000003_sig000001bf,
      LI => blk00000003_sig000001c0,
      O => blk00000003_sig000001c1
    );
  blk00000003_blk0000016f : XORCY
    port map (
      CI => blk00000003_sig000001bc,
      LI => blk00000003_sig000001bd,
      O => blk00000003_sig000001be
    );
  blk00000003_blk0000016e : XORCY
    port map (
      CI => blk00000003_sig000001bb,
      LI => NlwRenamedSig_OI_rfd,
      O => NLW_blk00000003_blk0000016e_O_UNCONNECTED
    );
  blk00000003_blk0000016d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(0),
      Q => blk00000003_sig000001ba
    );
  blk00000003_blk0000016c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(1),
      Q => blk00000003_sig000001b9
    );
  blk00000003_blk0000016b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(2),
      Q => blk00000003_sig000001b8
    );
  blk00000003_blk0000016a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(3),
      Q => blk00000003_sig000001b7
    );
  blk00000003_blk00000169 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(4),
      Q => blk00000003_sig000001b6
    );
  blk00000003_blk00000168 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(5),
      Q => blk00000003_sig000001b5
    );
  blk00000003_blk00000167 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(6),
      Q => blk00000003_sig000001b4
    );
  blk00000003_blk00000166 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(7),
      Q => blk00000003_sig000001b3
    );
  blk00000003_blk00000165 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(8),
      Q => blk00000003_sig000001b2
    );
  blk00000003_blk00000164 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(9),
      Q => blk00000003_sig000001b1
    );
  blk00000003_blk00000163 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(10),
      Q => blk00000003_sig000001b0
    );
  blk00000003_blk00000162 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(11),
      Q => blk00000003_sig000001af
    );
  blk00000003_blk00000161 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(12),
      Q => blk00000003_sig000001ae
    );
  blk00000003_blk00000160 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(13),
      Q => blk00000003_sig000001ad
    );
  blk00000003_blk0000015f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(14),
      Q => blk00000003_sig000001ac
    );
  blk00000003_blk0000015e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(15),
      Q => blk00000003_sig000001ab
    );
  blk00000003_blk0000015d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001ba,
      Q => blk00000003_sig000001aa
    );
  blk00000003_blk0000015c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001b9,
      Q => blk00000003_sig000001a9
    );
  blk00000003_blk0000015b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001b8,
      Q => blk00000003_sig000001a8
    );
  blk00000003_blk0000015a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001b7,
      Q => blk00000003_sig000001a7
    );
  blk00000003_blk00000159 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001b6,
      Q => blk00000003_sig000001a6
    );
  blk00000003_blk00000158 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001b5,
      Q => blk00000003_sig000001a5
    );
  blk00000003_blk00000157 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001b4,
      Q => blk00000003_sig000001a4
    );
  blk00000003_blk00000156 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001b3,
      Q => blk00000003_sig000001a3
    );
  blk00000003_blk00000155 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001b2,
      Q => blk00000003_sig000001a2
    );
  blk00000003_blk00000154 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001b1,
      Q => blk00000003_sig000001a1
    );
  blk00000003_blk00000153 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001b0,
      Q => blk00000003_sig000001a0
    );
  blk00000003_blk00000152 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001af,
      Q => blk00000003_sig0000019f
    );
  blk00000003_blk00000151 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001ae,
      Q => blk00000003_sig0000019e
    );
  blk00000003_blk00000150 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001ad,
      Q => blk00000003_sig0000019d
    );
  blk00000003_blk0000014f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001ac,
      Q => blk00000003_sig0000019c
    );
  blk00000003_blk0000014e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001ab,
      Q => blk00000003_sig0000019b
    );
  blk00000003_blk0000014d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001aa,
      Q => blk00000003_sig0000019a
    );
  blk00000003_blk0000014c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001a9,
      Q => blk00000003_sig00000199
    );
  blk00000003_blk0000014b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001a8,
      Q => blk00000003_sig00000198
    );
  blk00000003_blk0000014a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001a7,
      Q => blk00000003_sig00000197
    );
  blk00000003_blk00000149 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001a6,
      Q => blk00000003_sig00000196
    );
  blk00000003_blk00000148 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001a5,
      Q => blk00000003_sig00000195
    );
  blk00000003_blk00000147 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001a4,
      Q => blk00000003_sig00000194
    );
  blk00000003_blk00000146 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001a3,
      Q => blk00000003_sig00000193
    );
  blk00000003_blk00000145 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001a2,
      Q => blk00000003_sig00000192
    );
  blk00000003_blk00000144 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001a1,
      Q => blk00000003_sig00000191
    );
  blk00000003_blk00000143 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001a0,
      Q => blk00000003_sig00000190
    );
  blk00000003_blk00000142 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000019f,
      Q => blk00000003_sig0000018f
    );
  blk00000003_blk00000141 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000019e,
      Q => blk00000003_sig0000018e
    );
  blk00000003_blk00000140 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000019d,
      Q => blk00000003_sig0000018d
    );
  blk00000003_blk0000013f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000019c,
      Q => blk00000003_sig0000018c
    );
  blk00000003_blk0000013e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000019b,
      Q => blk00000003_sig0000018b
    );
  blk00000003_blk0000013d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000019a,
      Q => blk00000003_sig0000018a
    );
  blk00000003_blk0000013c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000199,
      Q => blk00000003_sig00000189
    );
  blk00000003_blk0000013b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000198,
      Q => blk00000003_sig00000188
    );
  blk00000003_blk0000013a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000197,
      Q => blk00000003_sig00000187
    );
  blk00000003_blk00000139 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000196,
      Q => blk00000003_sig00000186
    );
  blk00000003_blk00000138 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000195,
      Q => blk00000003_sig00000185
    );
  blk00000003_blk00000137 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000194,
      Q => blk00000003_sig00000184
    );
  blk00000003_blk00000136 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000193,
      Q => blk00000003_sig00000183
    );
  blk00000003_blk00000135 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000192,
      Q => blk00000003_sig00000182
    );
  blk00000003_blk00000134 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000191,
      Q => blk00000003_sig00000181
    );
  blk00000003_blk00000133 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000190,
      Q => blk00000003_sig00000180
    );
  blk00000003_blk00000132 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000018f,
      Q => blk00000003_sig0000017f
    );
  blk00000003_blk00000131 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000018e,
      Q => blk00000003_sig0000017e
    );
  blk00000003_blk00000130 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000018d,
      Q => blk00000003_sig0000017d
    );
  blk00000003_blk0000012f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000018c,
      Q => blk00000003_sig0000017c
    );
  blk00000003_blk0000012e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000018b,
      Q => blk00000003_sig0000017b
    );
  blk00000003_blk0000012d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000018a,
      Q => blk00000003_sig0000017a
    );
  blk00000003_blk0000012c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000189,
      Q => blk00000003_sig00000179
    );
  blk00000003_blk0000012b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000188,
      Q => blk00000003_sig00000178
    );
  blk00000003_blk0000012a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000187,
      Q => blk00000003_sig00000177
    );
  blk00000003_blk00000129 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000186,
      Q => blk00000003_sig00000176
    );
  blk00000003_blk00000128 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000185,
      Q => blk00000003_sig00000175
    );
  blk00000003_blk00000127 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000184,
      Q => blk00000003_sig00000174
    );
  blk00000003_blk00000126 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000183,
      Q => blk00000003_sig00000173
    );
  blk00000003_blk00000125 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000182,
      Q => blk00000003_sig00000172
    );
  blk00000003_blk00000124 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000181,
      Q => blk00000003_sig00000171
    );
  blk00000003_blk00000123 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000180,
      Q => blk00000003_sig00000170
    );
  blk00000003_blk00000122 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000017f,
      Q => blk00000003_sig0000016f
    );
  blk00000003_blk00000121 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000017e,
      Q => blk00000003_sig0000016e
    );
  blk00000003_blk00000120 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000017d,
      Q => blk00000003_sig0000016d
    );
  blk00000003_blk0000011f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000017c,
      Q => blk00000003_sig0000016c
    );
  blk00000003_blk0000011e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000017b,
      Q => blk00000003_sig0000016b
    );
  blk00000003_blk0000011d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000017a,
      Q => blk00000003_sig0000016a
    );
  blk00000003_blk0000011c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000179,
      Q => blk00000003_sig00000169
    );
  blk00000003_blk0000011b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000178,
      Q => blk00000003_sig00000168
    );
  blk00000003_blk0000011a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000177,
      Q => blk00000003_sig00000167
    );
  blk00000003_blk00000119 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000176,
      Q => blk00000003_sig00000166
    );
  blk00000003_blk00000118 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000175,
      Q => blk00000003_sig00000165
    );
  blk00000003_blk00000117 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000174,
      Q => blk00000003_sig00000164
    );
  blk00000003_blk00000116 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000173,
      Q => blk00000003_sig00000163
    );
  blk00000003_blk00000115 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000172,
      Q => blk00000003_sig00000162
    );
  blk00000003_blk00000114 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000171,
      Q => blk00000003_sig00000161
    );
  blk00000003_blk00000113 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000170,
      Q => blk00000003_sig00000160
    );
  blk00000003_blk00000112 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000016f,
      Q => blk00000003_sig0000015f
    );
  blk00000003_blk00000111 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000016e,
      Q => blk00000003_sig0000015e
    );
  blk00000003_blk00000110 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000016d,
      Q => blk00000003_sig0000015d
    );
  blk00000003_blk0000010f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000016c,
      Q => blk00000003_sig0000015c
    );
  blk00000003_blk0000010e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000016b,
      Q => blk00000003_sig0000015b
    );
  blk00000003_blk0000010d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000016a,
      Q => blk00000003_sig0000015a
    );
  blk00000003_blk0000010c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000169,
      Q => blk00000003_sig00000159
    );
  blk00000003_blk0000010b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000168,
      Q => blk00000003_sig00000158
    );
  blk00000003_blk0000010a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000167,
      Q => blk00000003_sig00000157
    );
  blk00000003_blk00000109 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000166,
      Q => blk00000003_sig00000156
    );
  blk00000003_blk00000108 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000165,
      Q => blk00000003_sig00000155
    );
  blk00000003_blk00000107 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000164,
      Q => blk00000003_sig00000154
    );
  blk00000003_blk00000106 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000163,
      Q => blk00000003_sig00000153
    );
  blk00000003_blk00000105 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000162,
      Q => blk00000003_sig00000152
    );
  blk00000003_blk00000104 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000161,
      Q => blk00000003_sig00000151
    );
  blk00000003_blk00000103 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000160,
      Q => blk00000003_sig00000150
    );
  blk00000003_blk00000102 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000015f,
      Q => blk00000003_sig0000014f
    );
  blk00000003_blk00000101 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000015e,
      Q => blk00000003_sig0000014e
    );
  blk00000003_blk00000100 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000015d,
      Q => blk00000003_sig0000014d
    );
  blk00000003_blk000000ff : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000015c,
      Q => blk00000003_sig0000014c
    );
  blk00000003_blk000000fe : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000015b,
      Q => blk00000003_sig0000014b
    );
  blk00000003_blk000000fd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000015a,
      Q => blk00000003_sig0000014a
    );
  blk00000003_blk000000fc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000159,
      Q => blk00000003_sig00000149
    );
  blk00000003_blk000000fb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000158,
      Q => blk00000003_sig00000148
    );
  blk00000003_blk000000fa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000157,
      Q => blk00000003_sig00000147
    );
  blk00000003_blk000000f9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000156,
      Q => blk00000003_sig00000146
    );
  blk00000003_blk000000f8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000155,
      Q => blk00000003_sig00000145
    );
  blk00000003_blk000000f7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000154,
      Q => blk00000003_sig00000144
    );
  blk00000003_blk000000f6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000153,
      Q => blk00000003_sig00000143
    );
  blk00000003_blk000000f5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000152,
      Q => blk00000003_sig00000142
    );
  blk00000003_blk000000f4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000151,
      Q => blk00000003_sig00000141
    );
  blk00000003_blk000000f3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000150,
      Q => blk00000003_sig00000140
    );
  blk00000003_blk000000f2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000014f,
      Q => blk00000003_sig0000013f
    );
  blk00000003_blk000000f1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000014e,
      Q => blk00000003_sig0000013e
    );
  blk00000003_blk000000f0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000014d,
      Q => blk00000003_sig0000013d
    );
  blk00000003_blk000000ef : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000014c,
      Q => blk00000003_sig0000013c
    );
  blk00000003_blk000000ee : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000014b,
      Q => blk00000003_sig0000013b
    );
  blk00000003_blk000000ed : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000014a,
      Q => blk00000003_sig0000013a
    );
  blk00000003_blk000000ec : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000149,
      Q => blk00000003_sig00000139
    );
  blk00000003_blk000000eb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000148,
      Q => blk00000003_sig00000138
    );
  blk00000003_blk000000ea : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000147,
      Q => blk00000003_sig00000137
    );
  blk00000003_blk000000e9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000146,
      Q => blk00000003_sig00000136
    );
  blk00000003_blk000000e8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000145,
      Q => blk00000003_sig00000135
    );
  blk00000003_blk000000e7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000144,
      Q => blk00000003_sig00000134
    );
  blk00000003_blk000000e6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000143,
      Q => blk00000003_sig00000133
    );
  blk00000003_blk000000e5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000142,
      Q => blk00000003_sig00000132
    );
  blk00000003_blk000000e4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000141,
      Q => blk00000003_sig00000131
    );
  blk00000003_blk000000e3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000140,
      Q => blk00000003_sig00000130
    );
  blk00000003_blk000000e2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000013f,
      Q => blk00000003_sig0000012f
    );
  blk00000003_blk000000e1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000013e,
      Q => blk00000003_sig0000012e
    );
  blk00000003_blk000000e0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000013d,
      Q => blk00000003_sig0000012d
    );
  blk00000003_blk000000df : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000013c,
      Q => blk00000003_sig0000012c
    );
  blk00000003_blk000000de : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000013b,
      Q => blk00000003_sig0000012b
    );
  blk00000003_blk000000dd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000013a,
      Q => blk00000003_sig0000012a
    );
  blk00000003_blk000000dc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000139,
      Q => blk00000003_sig00000129
    );
  blk00000003_blk000000db : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000138,
      Q => blk00000003_sig00000128
    );
  blk00000003_blk000000da : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000137,
      Q => blk00000003_sig00000127
    );
  blk00000003_blk000000d9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000136,
      Q => blk00000003_sig00000126
    );
  blk00000003_blk000000d8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000135,
      Q => blk00000003_sig00000125
    );
  blk00000003_blk000000d7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000134,
      Q => blk00000003_sig00000124
    );
  blk00000003_blk000000d6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000133,
      Q => blk00000003_sig00000123
    );
  blk00000003_blk000000d5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000132,
      Q => blk00000003_sig00000122
    );
  blk00000003_blk000000d4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000131,
      Q => blk00000003_sig00000121
    );
  blk00000003_blk000000d3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000130,
      Q => blk00000003_sig00000120
    );
  blk00000003_blk000000d2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000012f,
      Q => blk00000003_sig0000011f
    );
  blk00000003_blk000000d1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000012e,
      Q => blk00000003_sig0000011e
    );
  blk00000003_blk000000d0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000012d,
      Q => blk00000003_sig0000011d
    );
  blk00000003_blk000000cf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000012c,
      Q => blk00000003_sig0000011c
    );
  blk00000003_blk000000ce : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000012b,
      Q => blk00000003_sig0000011b
    );
  blk00000003_blk000000cd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000012a,
      Q => blk00000003_sig0000011a
    );
  blk00000003_blk000000cc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000129,
      Q => blk00000003_sig00000119
    );
  blk00000003_blk000000cb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000128,
      Q => blk00000003_sig00000118
    );
  blk00000003_blk000000ca : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000127,
      Q => blk00000003_sig00000117
    );
  blk00000003_blk000000c9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000126,
      Q => blk00000003_sig00000116
    );
  blk00000003_blk000000c8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000125,
      Q => blk00000003_sig00000115
    );
  blk00000003_blk000000c7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000124,
      Q => blk00000003_sig00000114
    );
  blk00000003_blk000000c6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000123,
      Q => blk00000003_sig00000113
    );
  blk00000003_blk000000c5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000122,
      Q => blk00000003_sig00000112
    );
  blk00000003_blk000000c4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000121,
      Q => blk00000003_sig00000111
    );
  blk00000003_blk000000c3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000120,
      Q => blk00000003_sig00000110
    );
  blk00000003_blk000000c2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000011f,
      Q => blk00000003_sig0000010f
    );
  blk00000003_blk000000c1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000011e,
      Q => blk00000003_sig0000010e
    );
  blk00000003_blk000000c0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000011d,
      Q => blk00000003_sig0000010d
    );
  blk00000003_blk000000bf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000011c,
      Q => blk00000003_sig0000010c
    );
  blk00000003_blk000000be : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000011b,
      Q => blk00000003_sig0000010b
    );
  blk00000003_blk000000bd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000011a,
      Q => blk00000003_sig0000010a
    );
  blk00000003_blk000000bc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000119,
      Q => blk00000003_sig00000109
    );
  blk00000003_blk000000bb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000118,
      Q => blk00000003_sig00000108
    );
  blk00000003_blk000000ba : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000117,
      Q => blk00000003_sig00000107
    );
  blk00000003_blk000000b9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000116,
      Q => blk00000003_sig00000106
    );
  blk00000003_blk000000b8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000115,
      Q => blk00000003_sig00000105
    );
  blk00000003_blk000000b7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000114,
      Q => blk00000003_sig00000104
    );
  blk00000003_blk000000b6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000113,
      Q => blk00000003_sig00000103
    );
  blk00000003_blk000000b5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000112,
      Q => blk00000003_sig00000102
    );
  blk00000003_blk000000b4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000111,
      Q => blk00000003_sig00000101
    );
  blk00000003_blk000000b3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000110,
      Q => blk00000003_sig00000100
    );
  blk00000003_blk000000b2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000010f,
      Q => blk00000003_sig000000ff
    );
  blk00000003_blk000000b1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000010e,
      Q => blk00000003_sig000000fe
    );
  blk00000003_blk000000b0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000010d,
      Q => blk00000003_sig000000fd
    );
  blk00000003_blk000000af : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000010c,
      Q => blk00000003_sig000000fc
    );
  blk00000003_blk000000ae : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000010b,
      Q => blk00000003_sig000000fb
    );
  blk00000003_blk000000ad : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000010a,
      Q => blk00000003_sig000000fa
    );
  blk00000003_blk000000ac : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000109,
      Q => blk00000003_sig000000f9
    );
  blk00000003_blk000000ab : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000108,
      Q => blk00000003_sig000000f8
    );
  blk00000003_blk000000aa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000107,
      Q => blk00000003_sig000000f7
    );
  blk00000003_blk000000a9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000106,
      Q => blk00000003_sig000000f6
    );
  blk00000003_blk000000a8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000105,
      Q => blk00000003_sig000000f5
    );
  blk00000003_blk000000a7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000104,
      Q => blk00000003_sig000000f4
    );
  blk00000003_blk000000a6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000103,
      Q => blk00000003_sig000000f3
    );
  blk00000003_blk000000a5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000102,
      Q => blk00000003_sig000000f2
    );
  blk00000003_blk000000a4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000101,
      Q => blk00000003_sig000000f1
    );
  blk00000003_blk000000a3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000100,
      Q => blk00000003_sig000000f0
    );
  blk00000003_blk000000a2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ff,
      Q => blk00000003_sig000000ef
    );
  blk00000003_blk000000a1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000fe,
      Q => blk00000003_sig000000ee
    );
  blk00000003_blk000000a0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000fd,
      Q => blk00000003_sig000000ed
    );
  blk00000003_blk0000009f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000fc,
      Q => blk00000003_sig000000ec
    );
  blk00000003_blk0000009e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000fb,
      Q => blk00000003_sig000000eb
    );
  blk00000003_blk0000009d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000fa,
      Q => blk00000003_sig000000ea
    );
  blk00000003_blk0000009c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f9,
      Q => blk00000003_sig000000e9
    );
  blk00000003_blk0000009b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f8,
      Q => blk00000003_sig000000e8
    );
  blk00000003_blk0000009a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f7,
      Q => blk00000003_sig000000e7
    );
  blk00000003_blk00000099 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f6,
      Q => blk00000003_sig000000e6
    );
  blk00000003_blk00000098 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f5,
      Q => blk00000003_sig000000e5
    );
  blk00000003_blk00000097 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f4,
      Q => blk00000003_sig000000e4
    );
  blk00000003_blk00000096 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f3,
      Q => blk00000003_sig000000e3
    );
  blk00000003_blk00000095 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f2,
      Q => blk00000003_sig000000e2
    );
  blk00000003_blk00000094 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f1,
      Q => blk00000003_sig000000e1
    );
  blk00000003_blk00000093 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f0,
      Q => blk00000003_sig000000e0
    );
  blk00000003_blk00000092 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ef,
      Q => blk00000003_sig000000df
    );
  blk00000003_blk00000091 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ee,
      Q => blk00000003_sig000000de
    );
  blk00000003_blk00000090 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ed,
      Q => blk00000003_sig000000dd
    );
  blk00000003_blk0000008f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ec,
      Q => blk00000003_sig000000dc
    );
  blk00000003_blk0000008e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000eb,
      Q => blk00000003_sig000000db
    );
  blk00000003_blk0000008d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ea,
      Q => blk00000003_sig000000da
    );
  blk00000003_blk0000008c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e9,
      Q => blk00000003_sig000000d9
    );
  blk00000003_blk0000008b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e8,
      Q => blk00000003_sig000000d8
    );
  blk00000003_blk0000008a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e7,
      Q => blk00000003_sig000000d7
    );
  blk00000003_blk00000089 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e6,
      Q => blk00000003_sig000000d6
    );
  blk00000003_blk00000088 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e5,
      Q => blk00000003_sig000000d5
    );
  blk00000003_blk00000087 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e4,
      Q => blk00000003_sig000000d4
    );
  blk00000003_blk00000086 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e3,
      Q => blk00000003_sig000000d3
    );
  blk00000003_blk00000085 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e2,
      Q => blk00000003_sig000000d2
    );
  blk00000003_blk00000084 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e1,
      Q => blk00000003_sig000000d1
    );
  blk00000003_blk00000083 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e0,
      Q => blk00000003_sig000000d0
    );
  blk00000003_blk00000082 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000df,
      Q => blk00000003_sig000000cf
    );
  blk00000003_blk00000081 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000de,
      Q => blk00000003_sig000000ce
    );
  blk00000003_blk00000080 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000dd,
      Q => blk00000003_sig000000cd
    );
  blk00000003_blk0000007f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000dc,
      Q => blk00000003_sig000000cc
    );
  blk00000003_blk0000007e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000db,
      Q => blk00000003_sig000000cb
    );
  blk00000003_blk0000007d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000da,
      Q => blk00000003_sig000000c9
    );
  blk00000003_blk0000007c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d9,
      Q => blk00000003_sig000000c7
    );
  blk00000003_blk0000007b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d8,
      Q => blk00000003_sig000000c5
    );
  blk00000003_blk0000007a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d7,
      Q => blk00000003_sig000000c3
    );
  blk00000003_blk00000079 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d6,
      Q => blk00000003_sig000000c1
    );
  blk00000003_blk00000078 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d5,
      Q => blk00000003_sig000000bf
    );
  blk00000003_blk00000077 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d4,
      Q => blk00000003_sig000000bd
    );
  blk00000003_blk00000076 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d3,
      Q => blk00000003_sig000000bb
    );
  blk00000003_blk00000075 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d2,
      Q => blk00000003_sig000000b9
    );
  blk00000003_blk00000074 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d1,
      Q => blk00000003_sig000000b7
    );
  blk00000003_blk00000073 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d0,
      Q => blk00000003_sig000000b5
    );
  blk00000003_blk00000072 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000cf,
      Q => blk00000003_sig000000b3
    );
  blk00000003_blk00000071 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ce,
      Q => blk00000003_sig000000b1
    );
  blk00000003_blk00000070 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000cd,
      Q => blk00000003_sig000000af
    );
  blk00000003_blk0000006f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000cc,
      Q => blk00000003_sig000000ad
    );
  blk00000003_blk0000006e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000cb,
      Q => blk00000003_sig000000ab
    );
  blk00000003_blk0000006d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c9,
      Q => blk00000003_sig000000ca
    );
  blk00000003_blk0000006c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c7,
      Q => blk00000003_sig000000c8
    );
  blk00000003_blk0000006b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c5,
      Q => blk00000003_sig000000c6
    );
  blk00000003_blk0000006a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c3,
      Q => blk00000003_sig000000c4
    );
  blk00000003_blk00000069 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c1,
      Q => blk00000003_sig000000c2
    );
  blk00000003_blk00000068 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000bf,
      Q => blk00000003_sig000000c0
    );
  blk00000003_blk00000067 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000bd,
      Q => blk00000003_sig000000be
    );
  blk00000003_blk00000066 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000bb,
      Q => blk00000003_sig000000bc
    );
  blk00000003_blk00000065 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b9,
      Q => blk00000003_sig000000ba
    );
  blk00000003_blk00000064 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b7,
      Q => blk00000003_sig000000b8
    );
  blk00000003_blk00000063 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b5,
      Q => blk00000003_sig000000b6
    );
  blk00000003_blk00000062 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b3,
      Q => blk00000003_sig000000b4
    );
  blk00000003_blk00000061 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b1,
      Q => blk00000003_sig000000b2
    );
  blk00000003_blk00000060 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000af,
      Q => blk00000003_sig000000b0
    );
  blk00000003_blk0000005f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ad,
      Q => blk00000003_sig000000ae
    );
  blk00000003_blk0000005e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ab,
      Q => blk00000003_sig000000ac
    );
  blk00000003_blk0000005d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(0),
      Q => blk00000003_sig000000aa
    );
  blk00000003_blk0000005c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(1),
      Q => blk00000003_sig000000a9
    );
  blk00000003_blk0000005b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(2),
      Q => blk00000003_sig000000a8
    );
  blk00000003_blk0000005a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(3),
      Q => blk00000003_sig000000a7
    );
  blk00000003_blk00000059 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(4),
      Q => blk00000003_sig000000a6
    );
  blk00000003_blk00000058 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(5),
      Q => blk00000003_sig000000a5
    );
  blk00000003_blk00000057 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(6),
      Q => blk00000003_sig000000a4
    );
  blk00000003_blk00000056 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(7),
      Q => blk00000003_sig000000a3
    );
  blk00000003_blk00000055 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(8),
      Q => blk00000003_sig000000a2
    );
  blk00000003_blk00000054 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(9),
      Q => blk00000003_sig000000a1
    );
  blk00000003_blk00000053 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(10),
      Q => blk00000003_sig000000a0
    );
  blk00000003_blk00000052 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(11),
      Q => blk00000003_sig0000009f
    );
  blk00000003_blk00000051 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(12),
      Q => blk00000003_sig0000009e
    );
  blk00000003_blk00000050 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(13),
      Q => blk00000003_sig0000009d
    );
  blk00000003_blk0000004f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(14),
      Q => blk00000003_sig0000009c
    );
  blk00000003_blk0000004e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(15),
      Q => blk00000003_sig0000009b
    );
  blk00000003_blk0000004d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000009a,
      Q => quotient(0)
    );
  blk00000003_blk0000004c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000099,
      Q => quotient(1)
    );
  blk00000003_blk0000004b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000098,
      Q => quotient(2)
    );
  blk00000003_blk0000004a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000097,
      Q => quotient(3)
    );
  blk00000003_blk00000049 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000096,
      Q => quotient(4)
    );
  blk00000003_blk00000048 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000095,
      Q => quotient(5)
    );
  blk00000003_blk00000047 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000094,
      Q => quotient(6)
    );
  blk00000003_blk00000046 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000093,
      Q => quotient(7)
    );
  blk00000003_blk00000045 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000092,
      Q => quotient(8)
    );
  blk00000003_blk00000044 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000091,
      Q => quotient(9)
    );
  blk00000003_blk00000043 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000090,
      Q => quotient(10)
    );
  blk00000003_blk00000042 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000008f,
      Q => quotient(11)
    );
  blk00000003_blk00000041 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000008e,
      Q => quotient(12)
    );
  blk00000003_blk00000040 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000008d,
      Q => quotient(13)
    );
  blk00000003_blk0000003f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000008c,
      Q => quotient(14)
    );
  blk00000003_blk0000003e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000008b,
      Q => quotient(15)
    );
  blk00000003_blk0000003d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000046,
      Q => blk00000003_sig0000008a
    );
  blk00000003_blk0000003c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000089,
      Q => blk00000003_sig00000088
    );
  blk00000003_blk0000003b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000088,
      Q => blk00000003_sig00000086
    );
  blk00000003_blk0000003a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000087,
      Q => blk00000003_sig00000085
    );
  blk00000003_blk00000039 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000086,
      Q => blk00000003_sig00000083
    );
  blk00000003_blk00000038 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000085,
      Q => blk00000003_sig00000082
    );
  blk00000003_blk00000037 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000084,
      Q => blk00000003_sig00000081
    );
  blk00000003_blk00000036 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000083,
      Q => blk00000003_sig0000007f
    );
  blk00000003_blk00000035 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000082,
      Q => blk00000003_sig0000007e
    );
  blk00000003_blk00000034 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000081,
      Q => blk00000003_sig0000007d
    );
  blk00000003_blk00000033 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000080,
      Q => blk00000003_sig0000007c
    );
  blk00000003_blk00000032 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007f,
      Q => blk00000003_sig0000007a
    );
  blk00000003_blk00000031 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007e,
      Q => blk00000003_sig00000079
    );
  blk00000003_blk00000030 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007d,
      Q => blk00000003_sig00000078
    );
  blk00000003_blk0000002f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007c,
      Q => blk00000003_sig00000077
    );
  blk00000003_blk0000002e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007b,
      Q => blk00000003_sig00000076
    );
  blk00000003_blk0000002d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007a,
      Q => blk00000003_sig00000073
    );
  blk00000003_blk0000002c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000079,
      Q => blk00000003_sig00000071
    );
  blk00000003_blk0000002b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000078,
      Q => blk00000003_sig0000006f
    );
  blk00000003_blk0000002a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000077,
      Q => blk00000003_sig0000006d
    );
  blk00000003_blk00000029 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000076,
      Q => blk00000003_sig0000006b
    );
  blk00000003_blk00000028 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000075,
      Q => blk00000003_sig00000069
    );
  blk00000003_blk00000027 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000073,
      Q => blk00000003_sig00000074
    );
  blk00000003_blk00000026 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000071,
      Q => blk00000003_sig00000072
    );
  blk00000003_blk00000025 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006f,
      Q => blk00000003_sig00000070
    );
  blk00000003_blk00000024 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006d,
      Q => blk00000003_sig0000006e
    );
  blk00000003_blk00000023 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006b,
      Q => blk00000003_sig0000006c
    );
  blk00000003_blk00000022 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000069,
      Q => blk00000003_sig0000006a
    );
  blk00000003_blk00000021 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000067,
      Q => blk00000003_sig00000068
    );
  blk00000003_blk00000020 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000065,
      Q => blk00000003_sig00000066
    );
  blk00000003_blk0000001f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000064,
      Q => blk00000003_sig0000005d
    );
  blk00000003_blk0000001e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000063,
      Q => blk00000003_sig0000005c
    );
  blk00000003_blk0000001d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000062,
      Q => blk00000003_sig0000005b
    );
  blk00000003_blk0000001c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000061,
      Q => blk00000003_sig0000005a
    );
  blk00000003_blk0000001b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000060,
      Q => blk00000003_sig00000059
    );
  blk00000003_blk0000001a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000005f,
      Q => blk00000003_sig00000058
    );
  blk00000003_blk00000019 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000005d,
      Q => blk00000003_sig0000005e
    );
  blk00000003_blk00000018 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000005c,
      Q => blk00000003_sig00000056
    );
  blk00000003_blk00000017 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000005b,
      Q => blk00000003_sig00000055
    );
  blk00000003_blk00000016 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000005a,
      Q => blk00000003_sig00000054
    );
  blk00000003_blk00000015 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000059,
      Q => blk00000003_sig00000053
    );
  blk00000003_blk00000014 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000058,
      Q => blk00000003_sig00000052
    );
  blk00000003_blk00000013 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000056,
      Q => blk00000003_sig00000057
    );
  blk00000003_blk00000012 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000055,
      Q => blk00000003_sig00000050
    );
  blk00000003_blk00000011 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000054,
      Q => blk00000003_sig0000004f
    );
  blk00000003_blk00000010 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000053,
      Q => blk00000003_sig0000004e
    );
  blk00000003_blk0000000f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000052,
      Q => blk00000003_sig0000004d
    );
  blk00000003_blk0000000e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000050,
      Q => blk00000003_sig00000051
    );
  blk00000003_blk0000000d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000004f,
      Q => blk00000003_sig0000004b
    );
  blk00000003_blk0000000c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000004e,
      Q => blk00000003_sig0000004a
    );
  blk00000003_blk0000000b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000004d,
      Q => blk00000003_sig00000049
    );
  blk00000003_blk0000000a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000004b,
      Q => blk00000003_sig0000004c
    );
  blk00000003_blk00000009 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000004a,
      Q => blk00000003_sig00000047
    );
  blk00000003_blk00000008 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000049,
      Q => blk00000003_sig00000045
    );
  blk00000003_blk00000007 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000047,
      Q => blk00000003_sig00000048
    );
  blk00000003_blk00000006 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000045,
      Q => blk00000003_sig00000046
    );
  blk00000003_blk00000005 : VCC
    port map (
      P => NlwRenamedSig_OI_rfd
    );
  blk00000003_blk00000004 : GND
    port map (
      G => blk00000003_sig00000043
    );

end STRUCTURE;

-- synthesis translate_on

-------------------------------------------------------------------
-- System Generator version 13.2 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
package conv_pkg is
    constant simulating : boolean := false
      -- synopsys translate_off
        or true
      -- synopsys translate_on
    ;
    constant xlUnsigned : integer := 1;
    constant xlSigned : integer := 2;
    constant xlWrap : integer := 1;
    constant xlSaturate : integer := 2;
    constant xlTruncate : integer := 1;
    constant xlRound : integer := 2;
    constant xlRoundBanker : integer := 3;
    constant xlAddMode : integer := 1;
    constant xlSubMode : integer := 2;
    attribute black_box : boolean;
    attribute syn_black_box : boolean;
    attribute fpga_dont_touch: string;
    attribute box_type :  string;
    attribute keep : string;
    attribute syn_keep : boolean;
    function std_logic_vector_to_unsigned(inp : std_logic_vector) return unsigned;
    function unsigned_to_std_logic_vector(inp : unsigned) return std_logic_vector;
    function std_logic_vector_to_signed(inp : std_logic_vector) return signed;
    function signed_to_std_logic_vector(inp : signed) return std_logic_vector;
    function unsigned_to_signed(inp : unsigned) return signed;
    function signed_to_unsigned(inp : signed) return unsigned;
    function pos(inp : std_logic_vector; arith : INTEGER) return boolean;
    function all_same(inp: std_logic_vector) return boolean;
    function all_zeros(inp: std_logic_vector) return boolean;
    function is_point_five(inp: std_logic_vector) return boolean;
    function all_ones(inp: std_logic_vector) return boolean;
    function convert_type (inp : std_logic_vector; old_width, old_bin_pt,
                           old_arith, new_width, new_bin_pt, new_arith,
                           quantization, overflow : INTEGER)
        return std_logic_vector;
    function cast (inp : std_logic_vector; old_bin_pt,
                   new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector;
    function vec_slice (inp : std_logic_vector; upper, lower : INTEGER)
        return std_logic_vector;
    function s2u_slice (inp : signed; upper, lower : INTEGER)
        return unsigned;
    function u2u_slice (inp : unsigned; upper, lower : INTEGER)
        return unsigned;
    function s2s_cast (inp : signed; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return signed;
    function u2s_cast (inp : unsigned; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return signed;
    function s2u_cast (inp : signed; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return unsigned;
    function u2u_cast (inp : unsigned; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return unsigned;
    function u2v_cast (inp : unsigned; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return std_logic_vector;
    function s2v_cast (inp : signed; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return std_logic_vector;
    function trunc (inp : std_logic_vector; old_width, old_bin_pt, old_arith,
                    new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector;
    function round_towards_inf (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt,
                                new_arith : INTEGER) return std_logic_vector;
    function round_towards_even (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt,
                                new_arith : INTEGER) return std_logic_vector;
    function max_signed(width : INTEGER) return std_logic_vector;
    function min_signed(width : INTEGER) return std_logic_vector;
    function saturation_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                              old_arith, new_width, new_bin_pt, new_arith
                              : INTEGER) return std_logic_vector;
    function wrap_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                        old_arith, new_width, new_bin_pt, new_arith : INTEGER)
                        return std_logic_vector;
    function fractional_bits(a_bin_pt, b_bin_pt: INTEGER) return INTEGER;
    function integer_bits(a_width, a_bin_pt, b_width, b_bin_pt: INTEGER)
        return INTEGER;
    function sign_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector;
    function zero_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector;
    function zero_ext(inp : std_logic; new_width : INTEGER)
        return std_logic_vector;
    function extend_MSB(inp : std_logic_vector; new_width, arith : INTEGER)
        return std_logic_vector;
    function align_input(inp : std_logic_vector; old_width, delta, new_arith,
                          new_width: INTEGER)
        return std_logic_vector;
    function pad_LSB(inp : std_logic_vector; new_width: integer)
        return std_logic_vector;
    function pad_LSB(inp : std_logic_vector; new_width, arith : integer)
        return std_logic_vector;
    function max(L, R: INTEGER) return INTEGER;
    function min(L, R: INTEGER) return INTEGER;
    function "="(left,right: STRING) return boolean;
    function boolean_to_signed (inp : boolean; width: integer)
        return signed;
    function boolean_to_unsigned (inp : boolean; width: integer)
        return unsigned;
    function boolean_to_vector (inp : boolean)
        return std_logic_vector;
    function std_logic_to_vector (inp : std_logic)
        return std_logic_vector;
    function integer_to_std_logic_vector (inp : integer;  width, arith : integer)
        return std_logic_vector;
    function std_logic_vector_to_integer (inp : std_logic_vector;  arith : integer)
        return integer;
    function std_logic_to_integer(constant inp : std_logic := '0')
        return integer;
    function bin_string_element_to_std_logic_vector (inp : string;  width, index : integer)
        return std_logic_vector;
    function bin_string_to_std_logic_vector (inp : string)
        return std_logic_vector;
    function hex_string_to_std_logic_vector (inp : string; width : integer)
        return std_logic_vector;
    function makeZeroBinStr (width : integer) return STRING;
    function and_reduce(inp: std_logic_vector) return std_logic;
    -- synopsys translate_off
    function is_binary_string_invalid (inp : string)
        return boolean;
    function is_binary_string_undefined (inp : string)
        return boolean;
    function is_XorU(inp : std_logic_vector)
        return boolean;
    function to_real(inp : std_logic_vector; bin_pt : integer; arith : integer)
        return real;
    function std_logic_to_real(inp : std_logic; bin_pt : integer; arith : integer)
        return real;
    function real_to_std_logic_vector (inp : real;  width, bin_pt, arith : integer)
        return std_logic_vector;
    function real_string_to_std_logic_vector (inp : string;  width, bin_pt, arith : integer)
        return std_logic_vector;
    constant display_precision : integer := 20;
    function real_to_string (inp : real) return string;
    function valid_bin_string(inp : string) return boolean;
    function std_logic_vector_to_bin_string(inp : std_logic_vector) return string;
    function std_logic_to_bin_string(inp : std_logic) return string;
    function std_logic_vector_to_bin_string_w_point(inp : std_logic_vector; bin_pt : integer)
        return string;
    function real_to_bin_string(inp : real;  width, bin_pt, arith : integer)
        return string;
    type stdlogic_to_char_t is array(std_logic) of character;
    constant to_char : stdlogic_to_char_t := (
        'U' => 'U',
        'X' => 'X',
        '0' => '0',
        '1' => '1',
        'Z' => 'Z',
        'W' => 'W',
        'L' => 'L',
        'H' => 'H',
        '-' => '-');
    -- synopsys translate_on
end conv_pkg;
package body conv_pkg is
    function std_logic_vector_to_unsigned(inp : std_logic_vector)
        return unsigned
    is
    begin
        return unsigned (inp);
    end;
    function unsigned_to_std_logic_vector(inp : unsigned)
        return std_logic_vector
    is
    begin
        return std_logic_vector(inp);
    end;
    function std_logic_vector_to_signed(inp : std_logic_vector)
        return signed
    is
    begin
        return  signed (inp);
    end;
    function signed_to_std_logic_vector(inp : signed)
        return std_logic_vector
    is
    begin
        return std_logic_vector(inp);
    end;
    function unsigned_to_signed (inp : unsigned)
        return signed
    is
    begin
        return signed(std_logic_vector(inp));
    end;
    function signed_to_unsigned (inp : signed)
        return unsigned
    is
    begin
        return unsigned(std_logic_vector(inp));
    end;
    function pos(inp : std_logic_vector; arith : INTEGER)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        if arith = xlUnsigned then
            return true;
        else
            if vec(width-1) = '0' then
                return true;
            else
                return false;
            end if;
        end if;
        return true;
    end;
    function max_signed(width : INTEGER)
        return std_logic_vector
    is
        variable ones : std_logic_vector(width-2 downto 0);
        variable result : std_logic_vector(width-1 downto 0);
    begin
        ones := (others => '1');
        result(width-1) := '0';
        result(width-2 downto 0) := ones;
        return result;
    end;
    function min_signed(width : INTEGER)
        return std_logic_vector
    is
        variable zeros : std_logic_vector(width-2 downto 0);
        variable result : std_logic_vector(width-1 downto 0);
    begin
        zeros := (others => '0');
        result(width-1) := '1';
        result(width-2 downto 0) := zeros;
        return result;
    end;
    function and_reduce(inp: std_logic_vector) return std_logic
    is
        variable result: std_logic;
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        result := vec(0);
        if width > 1 then
            for i in 1 to width-1 loop
                result := result and vec(i);
            end loop;
        end if;
        return result;
    end;
    function all_same(inp: std_logic_vector) return boolean
    is
        variable result: boolean;
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        result := true;
        if width > 0 then
            for i in 1 to width-1 loop
                if vec(i) /= vec(0) then
                    result := false;
                end if;
            end loop;
        end if;
        return result;
    end;
    function all_zeros(inp: std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable zero : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        zero := (others => '0');
        vec := inp;
        -- synopsys translate_off
        if (is_XorU(vec)) then
            return false;
        end if;
         -- synopsys translate_on
        if (std_logic_vector_to_unsigned(vec) = std_logic_vector_to_unsigned(zero)) then
            result := true;
        else
            result := false;
        end if;
        return result;
    end;
    function is_point_five(inp: std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        vec := inp;
        -- synopsys translate_off
        if (is_XorU(vec)) then
            return false;
        end if;
         -- synopsys translate_on
        if (width > 1) then
           if ((vec(width-1) = '1') and (all_zeros(vec(width-2 downto 0)) = true)) then
               result := true;
           else
               result := false;
           end if;
        else
           if (vec(width-1) = '1') then
               result := true;
           else
               result := false;
           end if;
        end if;
        return result;
    end;
    function all_ones(inp: std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable one : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        one := (others => '1');
        vec := inp;
        -- synopsys translate_off
        if (is_XorU(vec)) then
            return false;
        end if;
         -- synopsys translate_on
        if (std_logic_vector_to_unsigned(vec) = std_logic_vector_to_unsigned(one)) then
            result := true;
        else
            result := false;
        end if;
        return result;
    end;
    function full_precision_num_width(quantization, overflow, old_width,
                                      old_bin_pt, old_arith,
                                      new_width, new_bin_pt, new_arith : INTEGER)
        return integer
    is
        variable result : integer;
    begin
        result := old_width + 2;
        return result;
    end;
    function quantized_num_width(quantization, overflow, old_width, old_bin_pt,
                                 old_arith, new_width, new_bin_pt, new_arith
                                 : INTEGER)
        return integer
    is
        variable right_of_dp, left_of_dp, result : integer;
    begin
        right_of_dp := max(new_bin_pt, old_bin_pt);
        left_of_dp := max((new_width - new_bin_pt), (old_width - old_bin_pt));
        result := (old_width + 2) + (new_bin_pt - old_bin_pt);
        return result;
    end;
    function convert_type (inp : std_logic_vector; old_width, old_bin_pt,
                           old_arith, new_width, new_bin_pt, new_arith,
                           quantization, overflow : INTEGER)
        return std_logic_vector
    is
        constant fp_width : integer :=
            full_precision_num_width(quantization, overflow, old_width,
                                     old_bin_pt, old_arith, new_width,
                                     new_bin_pt, new_arith);
        constant fp_bin_pt : integer := old_bin_pt;
        constant fp_arith : integer := old_arith;
        variable full_precision_result : std_logic_vector(fp_width-1 downto 0);
        constant q_width : integer :=
            quantized_num_width(quantization, overflow, old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt, new_arith);
        constant q_bin_pt : integer := new_bin_pt;
        constant q_arith : integer := old_arith;
        variable quantized_result : std_logic_vector(q_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        result := (others => '0');
        full_precision_result := cast(inp, old_bin_pt, fp_width, fp_bin_pt,
                                      fp_arith);
        if (quantization = xlRound) then
            quantized_result := round_towards_inf(full_precision_result,
                                                  fp_width, fp_bin_pt,
                                                  fp_arith, q_width, q_bin_pt,
                                                  q_arith);
        elsif (quantization = xlRoundBanker) then
            quantized_result := round_towards_even(full_precision_result,
                                                  fp_width, fp_bin_pt,
                                                  fp_arith, q_width, q_bin_pt,
                                                  q_arith);
        else
            quantized_result := trunc(full_precision_result, fp_width, fp_bin_pt,
                                      fp_arith, q_width, q_bin_pt, q_arith);
        end if;
        if (overflow = xlSaturate) then
            result := saturation_arith(quantized_result, q_width, q_bin_pt,
                                       q_arith, new_width, new_bin_pt, new_arith);
        else
             result := wrap_arith(quantized_result, q_width, q_bin_pt, q_arith,
                                  new_width, new_bin_pt, new_arith);
        end if;
        return result;
    end;
    function cast (inp : std_logic_vector; old_bin_pt, new_width,
                   new_bin_pt, new_arith : INTEGER)
        return std_logic_vector
    is
        constant old_width : integer := inp'length;
        constant left_of_dp : integer := (new_width - new_bin_pt)
                                         - (old_width - old_bin_pt);
        constant right_of_dp : integer := (new_bin_pt - old_bin_pt);
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable j   : integer;
    begin
        vec := inp;
        for i in new_width-1 downto 0 loop
            j := i - right_of_dp;
            if ( j > old_width-1) then
                if (new_arith = xlUnsigned) then
                    result(i) := '0';
                else
                    result(i) := vec(old_width-1);
                end if;
            elsif ( j >= 0) then
                result(i) := vec(j);
            else
                result(i) := '0';
            end if;
        end loop;
        return result;
    end;
    function vec_slice (inp : std_logic_vector; upper, lower : INTEGER)
      return std_logic_vector
    is
    begin
        return inp(upper downto lower);
    end;
    function s2u_slice (inp : signed; upper, lower : INTEGER)
      return unsigned
    is
    begin
        return unsigned(vec_slice(std_logic_vector(inp), upper, lower));
    end;
    function u2u_slice (inp : unsigned; upper, lower : INTEGER)
      return unsigned
    is
    begin
        return unsigned(vec_slice(std_logic_vector(inp), upper, lower));
    end;
    function s2s_cast (inp : signed; old_bin_pt, new_width, new_bin_pt : INTEGER)
        return signed
    is
    begin
        return signed(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlSigned));
    end;
    function s2u_cast (inp : signed; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return unsigned
    is
    begin
        return unsigned(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlSigned));
    end;
    function u2s_cast (inp : unsigned; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return signed
    is
    begin
        return signed(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlUnsigned));
    end;
    function u2u_cast (inp : unsigned; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return unsigned
    is
    begin
        return unsigned(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlUnsigned));
    end;
    function u2v_cast (inp : unsigned; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return std_logic_vector
    is
    begin
        return cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlUnsigned);
    end;
    function s2v_cast (inp : signed; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return std_logic_vector
    is
    begin
        return cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlSigned);
    end;
    function boolean_to_signed (inp : boolean; width : integer)
        return signed
    is
        variable result : signed(width - 1 downto 0);
    begin
        result := (others => '0');
        if inp then
          result(0) := '1';
        else
          result(0) := '0';
        end if;
        return result;
    end;
    function boolean_to_unsigned (inp : boolean; width : integer)
        return unsigned
    is
        variable result : unsigned(width - 1 downto 0);
    begin
        result := (others => '0');
        if inp then
          result(0) := '1';
        else
          result(0) := '0';
        end if;
        return result;
    end;
    function boolean_to_vector (inp : boolean)
        return std_logic_vector
    is
        variable result : std_logic_vector(1 - 1 downto 0);
    begin
        result := (others => '0');
        if inp then
          result(0) := '1';
        else
          result(0) := '0';
        end if;
        return result;
    end;
    function std_logic_to_vector (inp : std_logic)
        return std_logic_vector
    is
        variable result : std_logic_vector(1 - 1 downto 0);
    begin
        result(0) := inp;
        return result;
    end;
    function trunc (inp : std_logic_vector; old_width, old_bin_pt, old_arith,
                                new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector
    is
        constant right_of_dp : integer := (old_bin_pt - new_bin_pt);
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if right_of_dp >= 0 then
            if new_arith = xlUnsigned then
                result := zero_ext(vec(old_width-1 downto right_of_dp), new_width);
            else
                result := sign_ext(vec(old_width-1 downto right_of_dp), new_width);
            end if;
        else
            if new_arith = xlUnsigned then
                result := zero_ext(pad_LSB(vec, old_width +
                                           abs(right_of_dp)), new_width);
            else
                result := sign_ext(pad_LSB(vec, old_width +
                                           abs(right_of_dp)), new_width);
            end if;
        end if;
        return result;
    end;
    function round_towards_inf (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt, new_arith
                                : INTEGER)
        return std_logic_vector
    is
        constant right_of_dp : integer := (old_bin_pt - new_bin_pt);
        constant expected_new_width : integer :=  old_width - right_of_dp  + 1;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable one_or_zero : std_logic_vector(new_width-1 downto 0);
        variable truncated_val : std_logic_vector(new_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if right_of_dp >= 0 then
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            else
                truncated_val := sign_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            end if;
        else
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            else
                truncated_val := sign_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            end if;
        end if;
        one_or_zero := (others => '0');
        if (new_arith = xlSigned) then
            if (vec(old_width-1) = '0') then
                one_or_zero(0) := '1';
            end if;
            if (right_of_dp >= 2) and (right_of_dp <= old_width) then
                if (all_zeros(vec(right_of_dp-2 downto 0)) = false) then
                    one_or_zero(0) := '1';
                end if;
            end if;
            if (right_of_dp >= 1) and (right_of_dp <= old_width) then
                if vec(right_of_dp-1) = '0' then
                    one_or_zero(0) := '0';
                end if;
            else
                one_or_zero(0) := '0';
            end if;
        else
            if (right_of_dp >= 1) and (right_of_dp <= old_width) then
                one_or_zero(0) :=  vec(right_of_dp-1);
            end if;
        end if;
        if new_arith = xlSigned then
            result := signed_to_std_logic_vector(std_logic_vector_to_signed(truncated_val) +
                                                 std_logic_vector_to_signed(one_or_zero));
        else
            result := unsigned_to_std_logic_vector(std_logic_vector_to_unsigned(truncated_val) +
                                                  std_logic_vector_to_unsigned(one_or_zero));
        end if;
        return result;
    end;
    function round_towards_even (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt, new_arith
                                : INTEGER)
        return std_logic_vector
    is
        constant right_of_dp : integer := (old_bin_pt - new_bin_pt);
        constant expected_new_width : integer :=  old_width - right_of_dp  + 1;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable one_or_zero : std_logic_vector(new_width-1 downto 0);
        variable truncated_val : std_logic_vector(new_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if right_of_dp >= 0 then
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            else
                truncated_val := sign_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            end if;
        else
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            else
                truncated_val := sign_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            end if;
        end if;
        one_or_zero := (others => '0');
        if (right_of_dp >= 1) and (right_of_dp <= old_width) then
            if (is_point_five(vec(right_of_dp-1 downto 0)) = false) then
                one_or_zero(0) :=  vec(right_of_dp-1);
            else
                one_or_zero(0) :=  vec(right_of_dp);
            end if;
        end if;
        if new_arith = xlSigned then
            result := signed_to_std_logic_vector(std_logic_vector_to_signed(truncated_val) +
                                                 std_logic_vector_to_signed(one_or_zero));
        else
            result := unsigned_to_std_logic_vector(std_logic_vector_to_unsigned(truncated_val) +
                                                  std_logic_vector_to_unsigned(one_or_zero));
        end if;
        return result;
    end;
    function saturation_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                              old_arith, new_width, new_bin_pt, new_arith
                              : INTEGER)
        return std_logic_vector
    is
        constant left_of_dp : integer := (old_width - old_bin_pt) -
                                         (new_width - new_bin_pt);
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable overflow : boolean;
    begin
        vec := inp;
        overflow := true;
        result := (others => '0');
        if (new_width >= old_width) then
            overflow := false;
        end if;
        if ((old_arith = xlSigned and new_arith = xlSigned) and (old_width > new_width)) then
            if all_same(vec(old_width-1 downto new_width-1)) then
                overflow := false;
            end if;
        end if;
        if (old_arith = xlSigned and new_arith = xlUnsigned) then
            if (old_width > new_width) then
                if all_zeros(vec(old_width-1 downto new_width)) then
                    overflow := false;
                end if;
            else
                if (old_width = new_width) then
                    if (vec(new_width-1) = '0') then
                        overflow := false;
                    end if;
                end if;
            end if;
        end if;
        if (old_arith = xlUnsigned and new_arith = xlUnsigned) then
            if (old_width > new_width) then
                if all_zeros(vec(old_width-1 downto new_width)) then
                    overflow := false;
                end if;
            else
                if (old_width = new_width) then
                    overflow := false;
                end if;
            end if;
        end if;
        if ((old_arith = xlUnsigned and new_arith = xlSigned) and (old_width > new_width)) then
            if all_same(vec(old_width-1 downto new_width-1)) then
                overflow := false;
            end if;
        end if;
        if overflow then
            if new_arith = xlSigned then
                if vec(old_width-1) = '0' then
                    result := max_signed(new_width);
                else
                    result := min_signed(new_width);
                end if;
            else
                if ((old_arith = xlSigned) and vec(old_width-1) = '1') then
                    result := (others => '0');
                else
                    result := (others => '1');
                end if;
            end if;
        else
            if (old_arith = xlSigned) and (new_arith = xlUnsigned) then
                if (vec(old_width-1) = '1') then
                    vec := (others => '0');
                end if;
            end if;
            if new_width <= old_width then
                result := vec(new_width-1 downto 0);
            else
                if new_arith = xlUnsigned then
                    result := zero_ext(vec, new_width);
                else
                    result := sign_ext(vec, new_width);
                end if;
            end if;
        end if;
        return result;
    end;
   function wrap_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                       old_arith, new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector
    is
        variable result : std_logic_vector(new_width-1 downto 0);
        variable result_arith : integer;
    begin
        if (old_arith = xlSigned) and (new_arith = xlUnsigned) then
            result_arith := xlSigned;
        end if;
        result := cast(inp, old_bin_pt, new_width, new_bin_pt, result_arith);
        return result;
    end;
    function fractional_bits(a_bin_pt, b_bin_pt: INTEGER) return INTEGER is
    begin
        return max(a_bin_pt, b_bin_pt);
    end;
    function integer_bits(a_width, a_bin_pt, b_width, b_bin_pt: INTEGER)
        return INTEGER is
    begin
        return  max(a_width - a_bin_pt, b_width - b_bin_pt);
    end;
    function pad_LSB(inp : std_logic_vector; new_width: integer)
        return STD_LOGIC_VECTOR
    is
        constant orig_width : integer := inp'length;
        variable vec : std_logic_vector(orig_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable pos : integer;
        constant pad_pos : integer := new_width - orig_width - 1;
    begin
        vec := inp;
        pos := new_width-1;
        if (new_width >= orig_width) then
            for i in orig_width-1 downto 0 loop
                result(pos) := vec(i);
                pos := pos - 1;
            end loop;
            if pad_pos >= 0 then
                for i in pad_pos downto 0 loop
                    result(i) := '0';
                end loop;
            end if;
        end if;
        return result;
    end;
    function sign_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector
    is
        constant old_width : integer := inp'length;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if new_width >= old_width then
            result(old_width-1 downto 0) := vec;
            if new_width-1 >= old_width then
                for i in new_width-1 downto old_width loop
                    result(i) := vec(old_width-1);
                end loop;
            end if;
        else
            result(new_width-1 downto 0) := vec(new_width-1 downto 0);
        end if;
        return result;
    end;
    function zero_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector
    is
        constant old_width : integer := inp'length;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if new_width >= old_width then
            result(old_width-1 downto 0) := vec;
            if new_width-1 >= old_width then
                for i in new_width-1 downto old_width loop
                    result(i) := '0';
                end loop;
            end if;
        else
            result(new_width-1 downto 0) := vec(new_width-1 downto 0);
        end if;
        return result;
    end;
    function zero_ext(inp : std_logic; new_width : INTEGER)
        return std_logic_vector
    is
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        result(0) := inp;
        for i in new_width-1 downto 1 loop
            result(i) := '0';
        end loop;
        return result;
    end;
    function extend_MSB(inp : std_logic_vector; new_width, arith : INTEGER)
        return std_logic_vector
    is
        constant orig_width : integer := inp'length;
        variable vec : std_logic_vector(orig_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if arith = xlUnsigned then
            result := zero_ext(vec, new_width);
        else
            result := sign_ext(vec, new_width);
        end if;
        return result;
    end;
    function pad_LSB(inp : std_logic_vector; new_width, arith: integer)
        return STD_LOGIC_VECTOR
    is
        constant orig_width : integer := inp'length;
        variable vec : std_logic_vector(orig_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable pos : integer;
    begin
        vec := inp;
        pos := new_width-1;
        if (arith = xlUnsigned) then
            result(pos) := '0';
            pos := pos - 1;
        else
            result(pos) := vec(orig_width-1);
            pos := pos - 1;
        end if;
        if (new_width >= orig_width) then
            for i in orig_width-1 downto 0 loop
                result(pos) := vec(i);
                pos := pos - 1;
            end loop;
            if pos >= 0 then
                for i in pos downto 0 loop
                    result(i) := '0';
                end loop;
            end if;
        end if;
        return result;
    end;
    function align_input(inp : std_logic_vector; old_width, delta, new_arith,
                         new_width: INTEGER)
        return std_logic_vector
    is
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable padded_inp : std_logic_vector((old_width + delta)-1  downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if delta > 0 then
            padded_inp := pad_LSB(vec, old_width+delta);
            result := extend_MSB(padded_inp, new_width, new_arith);
        else
            result := extend_MSB(vec, new_width, new_arith);
        end if;
        return result;
    end;
    function max(L, R: INTEGER) return INTEGER is
    begin
        if L > R then
            return L;
        else
            return R;
        end if;
    end;
    function min(L, R: INTEGER) return INTEGER is
    begin
        if L < R then
            return L;
        else
            return R;
        end if;
    end;
    function "="(left,right: STRING) return boolean is
    begin
        if (left'length /= right'length) then
            return false;
        else
            test : for i in 1 to left'length loop
                if left(i) /= right(i) then
                    return false;
                end if;
            end loop test;
            return true;
        end if;
    end;
    -- synopsys translate_off
    function is_binary_string_invalid (inp : string)
        return boolean
    is
        variable vec : string(1 to inp'length);
        variable result : boolean;
    begin
        vec := inp;
        result := false;
        for i in 1 to vec'length loop
            if ( vec(i) = 'X' ) then
                result := true;
            end if;
        end loop;
        return result;
    end;
    function is_binary_string_undefined (inp : string)
        return boolean
    is
        variable vec : string(1 to inp'length);
        variable result : boolean;
    begin
        vec := inp;
        result := false;
        for i in 1 to vec'length loop
            if ( vec(i) = 'U' ) then
                result := true;
            end if;
        end loop;
        return result;
    end;
    function is_XorU(inp : std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        vec := inp;
        result := false;
        for i in 0 to width-1 loop
            if (vec(i) = 'U') or (vec(i) = 'X') then
                result := true;
            end if;
        end loop;
        return result;
    end;
    function to_real(inp : std_logic_vector; bin_pt : integer; arith : integer)
        return real
    is
        variable  vec : std_logic_vector(inp'length-1 downto 0);
        variable result, shift_val, undefined_real : real;
        variable neg_num : boolean;
    begin
        vec := inp;
        result := 0.0;
        neg_num := false;
        if vec(inp'length-1) = '1' then
            neg_num := true;
        end if;
        for i in 0 to inp'length-1 loop
            if  vec(i) = 'U' or vec(i) = 'X' then
                return undefined_real;
            end if;
            if arith = xlSigned then
                if neg_num then
                    if vec(i) = '0' then
                        result := result + 2.0**i;
                    end if;
                else
                    if vec(i) = '1' then
                        result := result + 2.0**i;
                    end if;
                end if;
            else
                if vec(i) = '1' then
                    result := result + 2.0**i;
                end if;
            end if;
        end loop;
        if arith = xlSigned then
            if neg_num then
                result := result + 1.0;
                result := result * (-1.0);
            end if;
        end if;
        shift_val := 2.0**(-1*bin_pt);
        result := result * shift_val;
        return result;
    end;
    function std_logic_to_real(inp : std_logic; bin_pt : integer; arith : integer)
        return real
    is
        variable result : real := 0.0;
    begin
        if inp = '1' then
            result := 1.0;
        end if;
        if arith = xlSigned then
            assert false
                report "It doesn't make sense to convert a 1 bit number to a signed real.";
        end if;
        return result;
    end;
    -- synopsys translate_on
    function integer_to_std_logic_vector (inp : integer;  width, arith : integer)
        return std_logic_vector
    is
        variable result : std_logic_vector(width-1 downto 0);
        variable unsigned_val : unsigned(width-1 downto 0);
        variable signed_val : signed(width-1 downto 0);
    begin
        if (arith = xlSigned) then
            signed_val := to_signed(inp, width);
            result := signed_to_std_logic_vector(signed_val);
        else
            unsigned_val := to_unsigned(inp, width);
            result := unsigned_to_std_logic_vector(unsigned_val);
        end if;
        return result;
    end;
    function std_logic_vector_to_integer (inp : std_logic_vector;  arith : integer)
        return integer
    is
        constant width : integer := inp'length;
        variable unsigned_val : unsigned(width-1 downto 0);
        variable signed_val : signed(width-1 downto 0);
        variable result : integer;
    begin
        if (arith = xlSigned) then
            signed_val := std_logic_vector_to_signed(inp);
            result := to_integer(signed_val);
        else
            unsigned_val := std_logic_vector_to_unsigned(inp);
            result := to_integer(unsigned_val);
        end if;
        return result;
    end;
    function std_logic_to_integer(constant inp : std_logic := '0')
        return integer
    is
    begin
        if inp = '1' then
            return 1;
        else
            return 0;
        end if;
    end;
    function makeZeroBinStr (width : integer) return STRING is
        variable result : string(1 to width+3);
    begin
        result(1) := '0';
        result(2) := 'b';
        for i in 3 to width+2 loop
            result(i) := '0';
        end loop;
        result(width+3) := '.';
        return result;
    end;
    -- synopsys translate_off
    function real_string_to_std_logic_vector (inp : string;  width, bin_pt, arith : integer)
        return std_logic_vector
    is
        variable result : std_logic_vector(width-1 downto 0);
    begin
        result := (others => '0');
        return result;
    end;
    function real_to_std_logic_vector (inp : real;  width, bin_pt, arith : integer)
        return std_logic_vector
    is
        variable real_val : real;
        variable int_val : integer;
        variable result : std_logic_vector(width-1 downto 0) := (others => '0');
        variable unsigned_val : unsigned(width-1 downto 0) := (others => '0');
        variable signed_val : signed(width-1 downto 0) := (others => '0');
    begin
        real_val := inp;
        int_val := integer(real_val * 2.0**(bin_pt));
        if (arith = xlSigned) then
            signed_val := to_signed(int_val, width);
            result := signed_to_std_logic_vector(signed_val);
        else
            unsigned_val := to_unsigned(int_val, width);
            result := unsigned_to_std_logic_vector(unsigned_val);
        end if;
        return result;
    end;
    -- synopsys translate_on
    function valid_bin_string (inp : string)
        return boolean
    is
        variable vec : string(1 to inp'length);
    begin
        vec := inp;
        if (vec(1) = '0' and vec(2) = 'b') then
            return true;
        else
            return false;
        end if;
    end;
    function hex_string_to_std_logic_vector(inp: string; width : integer)
        return std_logic_vector is
        constant strlen       : integer := inp'LENGTH;
        variable result       : std_logic_vector(width-1 downto 0);
        variable bitval       : std_logic_vector((strlen*4)-1 downto 0);
        variable posn         : integer;
        variable ch           : character;
        variable vec          : string(1 to strlen);
    begin
        vec := inp;
        result := (others => '0');
        posn := (strlen*4)-1;
        for i in 1 to strlen loop
            ch := vec(i);
            case ch is
                when '0' => bitval(posn downto posn-3) := "0000";
                when '1' => bitval(posn downto posn-3) := "0001";
                when '2' => bitval(posn downto posn-3) := "0010";
                when '3' => bitval(posn downto posn-3) := "0011";
                when '4' => bitval(posn downto posn-3) := "0100";
                when '5' => bitval(posn downto posn-3) := "0101";
                when '6' => bitval(posn downto posn-3) := "0110";
                when '7' => bitval(posn downto posn-3) := "0111";
                when '8' => bitval(posn downto posn-3) := "1000";
                when '9' => bitval(posn downto posn-3) := "1001";
                when 'A' | 'a' => bitval(posn downto posn-3) := "1010";
                when 'B' | 'b' => bitval(posn downto posn-3) := "1011";
                when 'C' | 'c' => bitval(posn downto posn-3) := "1100";
                when 'D' | 'd' => bitval(posn downto posn-3) := "1101";
                when 'E' | 'e' => bitval(posn downto posn-3) := "1110";
                when 'F' | 'f' => bitval(posn downto posn-3) := "1111";
                when others => bitval(posn downto posn-3) := "XXXX";
                               -- synopsys translate_off
                               ASSERT false
                                   REPORT "Invalid hex value" SEVERITY ERROR;
                               -- synopsys translate_on
            end case;
            posn := posn - 4;
        end loop;
        if (width <= strlen*4) then
            result :=  bitval(width-1 downto 0);
        else
            result((strlen*4)-1 downto 0) := bitval;
        end if;
        return result;
    end;
    function bin_string_to_std_logic_vector (inp : string)
        return std_logic_vector
    is
        variable pos : integer;
        variable vec : string(1 to inp'length);
        variable result : std_logic_vector(inp'length-1 downto 0);
    begin
        vec := inp;
        pos := inp'length-1;
        result := (others => '0');
        for i in 1 to vec'length loop
            -- synopsys translate_off
            if (pos < 0) and (vec(i) = '0' or vec(i) = '1' or vec(i) = 'X' or vec(i) = 'U')  then
                assert false
                    report "Input string is larger than output std_logic_vector. Truncating output.";
                return result;
            end if;
            -- synopsys translate_on
            if vec(i) = '0' then
                result(pos) := '0';
                pos := pos - 1;
            end if;
            if vec(i) = '1' then
                result(pos) := '1';
                pos := pos - 1;
            end if;
            -- synopsys translate_off
            if (vec(i) = 'X' or vec(i) = 'U') then
                result(pos) := 'U';
                pos := pos - 1;
            end if;
            -- synopsys translate_on
        end loop;
        return result;
    end;
    function bin_string_element_to_std_logic_vector (inp : string;  width, index : integer)
        return std_logic_vector
    is
        constant str_width : integer := width + 4;
        constant inp_len : integer := inp'length;
        constant num_elements : integer := (inp_len + 1)/str_width;
        constant reverse_index : integer := (num_elements-1) - index;
        variable left_pos : integer;
        variable right_pos : integer;
        variable vec : string(1 to inp'length);
        variable result : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        result := (others => '0');
        if (reverse_index = 0) and (reverse_index < num_elements) and (inp_len-3 >= width) then
            left_pos := 1;
            right_pos := width + 3;
            result := bin_string_to_std_logic_vector(vec(left_pos to right_pos));
        end if;
        if (reverse_index > 0) and (reverse_index < num_elements) and (inp_len-3 >= width) then
            left_pos := (reverse_index * str_width) + 1;
            right_pos := left_pos + width + 2;
            result := bin_string_to_std_logic_vector(vec(left_pos to right_pos));
        end if;
        return result;
    end;
   -- synopsys translate_off
    function std_logic_vector_to_bin_string(inp : std_logic_vector)
        return string
    is
        variable vec : std_logic_vector(1 to inp'length);
        variable result : string(vec'range);
    begin
        vec := inp;
        for i in vec'range loop
            result(i) := to_char(vec(i));
        end loop;
        return result;
    end;
    function std_logic_to_bin_string(inp : std_logic)
        return string
    is
        variable result : string(1 to 3);
    begin
        result(1) := '0';
        result(2) := 'b';
        result(3) := to_char(inp);
        return result;
    end;
    function std_logic_vector_to_bin_string_w_point(inp : std_logic_vector; bin_pt : integer)
        return string
    is
        variable width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable str_pos : integer;
        variable result : string(1 to width+3);
    begin
        vec := inp;
        str_pos := 1;
        result(str_pos) := '0';
        str_pos := 2;
        result(str_pos) := 'b';
        str_pos := 3;
        for i in width-1 downto 0  loop
            if (((width+3) - bin_pt) = str_pos) then
                result(str_pos) := '.';
                str_pos := str_pos + 1;
            end if;
            result(str_pos) := to_char(vec(i));
            str_pos := str_pos + 1;
        end loop;
        if (bin_pt = 0) then
            result(str_pos) := '.';
        end if;
        return result;
    end;
    function real_to_bin_string(inp : real;  width, bin_pt, arith : integer)
        return string
    is
        variable result : string(1 to width);
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := real_to_std_logic_vector(inp, width, bin_pt, arith);
        result := std_logic_vector_to_bin_string(vec);
        return result;
    end;
    function real_to_string (inp : real) return string
    is
        variable result : string(1 to display_precision) := (others => ' ');
    begin
        result(real'image(inp)'range) := real'image(inp);
        return result;
    end;
    -- synopsys translate_on
end conv_pkg;

-------------------------------------------------------------------
-- System Generator version 13.2 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
library block_id_calc_lib;
use block_id_calc_lib.conv_pkg.all;
entity srl17e is
    generic (width : integer:=16;
             latency : integer :=8);
    port (clk   : in std_logic;
          ce    : in std_logic;
          d     : in std_logic_vector(width-1 downto 0);
          q     : out std_logic_vector(width-1 downto 0));
end srl17e;
architecture structural of srl17e is
    component SRL16E
        port (D   : in STD_ULOGIC;
              CE  : in STD_ULOGIC;
              CLK : in STD_ULOGIC;
              A0  : in STD_ULOGIC;
              A1  : in STD_ULOGIC;
              A2  : in STD_ULOGIC;
              A3  : in STD_ULOGIC;
              Q   : out STD_ULOGIC);
    end component;
    attribute syn_black_box of SRL16E : component is true;
    attribute fpga_dont_touch of SRL16E : component is "true";
    component FDE
        port(
            Q  :        out   STD_ULOGIC;
            D  :        in    STD_ULOGIC;
            C  :        in    STD_ULOGIC;
            CE :        in    STD_ULOGIC);
    end component;
    attribute syn_black_box of FDE : component is true;
    attribute fpga_dont_touch of FDE : component is "true";
    constant a : std_logic_vector(4 downto 0) :=
        integer_to_std_logic_vector(latency-2,5,xlSigned);
    signal d_delayed : std_logic_vector(width-1 downto 0);
    signal srl16_out : std_logic_vector(width-1 downto 0);
begin
    d_delayed <= d after 200 ps;
    reg_array : for i in 0 to width-1 generate
        srl16_used: if latency > 1 generate
            u1 : srl16e port map(clk => clk,
                                 d => d_delayed(i),
                                 q => srl16_out(i),
                                 ce => ce,
                                 a0 => a(0),
                                 a1 => a(1),
                                 a2 => a(2),
                                 a3 => a(3));
        end generate;
        srl16_not_used: if latency <= 1 generate
            srl16_out(i) <= d_delayed(i);
        end generate;
        fde_used: if latency /= 0  generate
            u2 : fde port map(c => clk,
                              d => srl16_out(i),
                              q => q(i),
                              ce => ce);
        end generate;
        fde_not_used: if latency = 0  generate
            q(i) <= srl16_out(i);
        end generate;
    end generate;
 end structural;
library IEEE;
use IEEE.std_logic_1164.all;
library block_id_calc_lib;
use block_id_calc_lib.conv_pkg.all;
entity synth_reg is
    generic (width           : integer := 8;
             latency         : integer := 1);
    port (i       : in std_logic_vector(width-1 downto 0);
          ce      : in std_logic;
          clr     : in std_logic;
          clk     : in std_logic;
          o       : out std_logic_vector(width-1 downto 0));
end synth_reg;
architecture structural of synth_reg is
    component srl17e
        generic (width : integer:=16;
                 latency : integer :=8);
        port (clk : in std_logic;
              ce  : in std_logic;
              d   : in std_logic_vector(width-1 downto 0);
              q   : out std_logic_vector(width-1 downto 0));
    end component;
    function calc_num_srl17es (latency : integer)
        return integer
    is
        variable remaining_latency : integer;
        variable result : integer;
    begin
        result := latency / 17;
        remaining_latency := latency - (result * 17);
        if (remaining_latency /= 0) then
            result := result + 1;
        end if;
        return result;
    end;
    constant complete_num_srl17es : integer := latency / 17;
    constant num_srl17es : integer := calc_num_srl17es(latency);
    constant remaining_latency : integer := latency - (complete_num_srl17es * 17);
    type register_array is array (num_srl17es downto 0) of
        std_logic_vector(width-1 downto 0);
    signal z : register_array;
begin
    z(0) <= i;
    complete_ones : if complete_num_srl17es > 0 generate
        srl17e_array: for i in 0 to complete_num_srl17es-1 generate
            delay_comp : srl17e
                generic map (width => width,
                             latency => 17)
                port map (clk => clk,
                          ce  => ce,
                          d       => z(i),
                          q       => z(i+1));
        end generate;
    end generate;
    partial_one : if remaining_latency > 0 generate
        last_srl17e : srl17e
            generic map (width => width,
                         latency => remaining_latency)
            port map (clk => clk,
                      ce  => ce,
                      d   => z(num_srl17es-1),
                      q   => z(num_srl17es));
    end generate;
    o <= z(num_srl17es);
end structural;
library IEEE;
use IEEE.std_logic_1164.all;
library block_id_calc_lib;
use block_id_calc_lib.conv_pkg.all;
entity synth_reg_reg is
    generic (width           : integer := 8;
             latency         : integer := 1);
    port (i       : in std_logic_vector(width-1 downto 0);
          ce      : in std_logic;
          clr     : in std_logic;
          clk     : in std_logic;
          o       : out std_logic_vector(width-1 downto 0));
end synth_reg_reg;
architecture behav of synth_reg_reg is
  type reg_array_type is array (latency-1 downto 0) of std_logic_vector(width -1 downto 0);
  signal reg_bank : reg_array_type := (others => (others => '0'));
  signal reg_bank_in : reg_array_type := (others => (others => '0'));
  attribute syn_allow_retiming : boolean;
  attribute syn_srlstyle : string;
  attribute syn_allow_retiming of reg_bank : signal is true;
  attribute syn_allow_retiming of reg_bank_in : signal is true;
  attribute syn_srlstyle of reg_bank : signal is "registers";
  attribute syn_srlstyle of reg_bank_in : signal is "registers";
begin
  latency_eq_0: if latency = 0 generate
    o <= i;
  end generate latency_eq_0;
  latency_gt_0: if latency >= 1 generate
    o <= reg_bank(latency-1);
    reg_bank_in(0) <= i;
    loop_gen: for idx in latency-2 downto 0 generate
      reg_bank_in(idx+1) <= reg_bank(idx);
    end generate loop_gen;
    sync_loop: for sync_idx in latency-1 downto 0 generate
      sync_proc: process (clk)
      begin
        if clk'event and clk = '1' then
          if ce = '1'  then
            reg_bank(sync_idx) <= reg_bank_in(sync_idx);
          end if;
        end if;
      end process sync_proc;
    end generate sync_loop;
  end generate latency_gt_0;
end behav;

-------------------------------------------------------------------
-- System Generator version 13.2 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
library block_id_calc_lib;
use block_id_calc_lib.conv_pkg.all;
entity single_reg_w_init is
  generic (
    width: integer := 8;
    init_index: integer := 0;
    init_value: bit_vector := b"0000"
  );
  port (
    i: in std_logic_vector(width - 1 downto 0);
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    o: out std_logic_vector(width - 1 downto 0)
  );
end single_reg_w_init;
architecture structural of single_reg_w_init is
  function build_init_const(width: integer;
                            init_index: integer;
                            init_value: bit_vector)
    return std_logic_vector
  is
    variable result: std_logic_vector(width - 1 downto 0);
  begin
    if init_index = 0 then
      result := (others => '0');
    elsif init_index = 1 then
      result := (others => '0');
      result(0) := '1';
    else
      result := to_stdlogicvector(init_value);
    end if;
    return result;
  end;
  component fdre
    port (
      q: out std_ulogic;
      d: in  std_ulogic;
      c: in  std_ulogic;
      ce: in  std_ulogic;
      r: in  std_ulogic
    );
  end component;
  attribute syn_black_box of fdre: component is true;
  attribute fpga_dont_touch of fdre: component is "true";
  component fdse
    port (
      q: out std_ulogic;
      d: in  std_ulogic;
      c: in  std_ulogic;
      ce: in  std_ulogic;
      s: in  std_ulogic
    );
  end component;
  attribute syn_black_box of fdse: component is true;
  attribute fpga_dont_touch of fdse: component is "true";
  constant init_const: std_logic_vector(width - 1 downto 0)
    := build_init_const(width, init_index, init_value);
begin
  fd_prim_array: for index in 0 to width - 1 generate
    bit_is_0: if (init_const(index) = '0') generate
      fdre_comp: fdre
        port map (
          c => clk,
          d => i(index),
          q => o(index),
          ce => ce,
          r => clr
        );
    end generate;
    bit_is_1: if (init_const(index) = '1') generate
      fdse_comp: fdse
        port map (
          c => clk,
          d => i(index),
          q => o(index),
          ce => ce,
          s => clr
        );
    end generate;
  end generate;
end architecture structural;
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
library block_id_calc_lib;
use block_id_calc_lib.conv_pkg.all;
entity synth_reg_w_init is
  generic (
    width: integer := 8;
    init_index: integer := 0;
    init_value: bit_vector := b"0000";
    latency: integer := 1
  );
  port (
    i: in std_logic_vector(width - 1 downto 0);
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    o: out std_logic_vector(width - 1 downto 0)
  );
end synth_reg_w_init;
architecture structural of synth_reg_w_init is
  component single_reg_w_init
    generic (
      width: integer := 8;
      init_index: integer := 0;
      init_value: bit_vector := b"0000"
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  signal dly_i: std_logic_vector((latency + 1) * width - 1 downto 0);
  signal dly_clr: std_logic;
begin
  latency_eq_0: if (latency = 0) generate
    o <= i;
  end generate;
  latency_gt_0: if (latency >= 1) generate
    dly_i((latency + 1) * width - 1 downto latency * width) <= i
      after 200 ps;
    dly_clr <= clr after 200 ps;
    fd_array: for index in latency downto 1 generate
       reg_comp: single_reg_w_init
          generic map (
            width => width,
            init_index => init_index,
            init_value => init_value
          )
          port map (
            clk => clk,
            i => dly_i((index + 1) * width - 1 downto index * width),
            o => dly_i(index * width - 1 downto (index - 1) * width),
            ce => ce,
            clr => dly_clr
          );
    end generate;
    o <= dly_i(width - 1 downto 0);
  end generate;
end structural;

-------------------------------------------------------------------
-- System Generator version 13.2 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
library block_id_calc_lib;
use block_id_calc_lib.conv_pkg.all;
entity xladdsub is
  generic (
    core_name0: string := "";
    a_width: integer := 16;
    a_bin_pt: integer := 4;
    a_arith: integer := xlUnsigned;
    c_in_width: integer := 16;
    c_in_bin_pt: integer := 4;
    c_in_arith: integer := xlUnsigned;
    c_out_width: integer := 16;
    c_out_bin_pt: integer := 4;
    c_out_arith: integer := xlUnsigned;
    b_width: integer := 8;
    b_bin_pt: integer := 2;
    b_arith: integer := xlUnsigned;
    s_width: integer := 17;
    s_bin_pt: integer := 4;
    s_arith: integer := xlUnsigned;
    rst_width: integer := 1;
    rst_bin_pt: integer := 0;
    rst_arith: integer := xlUnsigned;
    en_width: integer := 1;
    en_bin_pt: integer := 0;
    en_arith: integer := xlUnsigned;
    full_s_width: integer := 17;
    full_s_arith: integer := xlUnsigned;
    mode: integer := xlAddMode;
    extra_registers: integer := 0;
    latency: integer := 0;
    quantization: integer := xlTruncate;
    overflow: integer := xlWrap;
    c_latency: integer := 0;
    c_output_width: integer := 17;
    c_has_c_in : integer := 0;
    c_has_c_out : integer := 0
  );
  port (
    a: in std_logic_vector(a_width - 1 downto 0);
    b: in std_logic_vector(b_width - 1 downto 0);
    c_in : in std_logic_vector (0 downto 0) := "0";
    ce: in std_logic;
    clr: in std_logic := '0';
    clk: in std_logic;
    rst: in std_logic_vector(rst_width - 1 downto 0) := "0";
    en: in std_logic_vector(en_width - 1 downto 0) := "1";
    c_out : out std_logic_vector (0 downto 0);
    s: out std_logic_vector(s_width - 1 downto 0)
  );
end xladdsub;
architecture behavior of xladdsub is
  component synth_reg
    generic (
      width: integer := 16;
      latency: integer := 5
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  function format_input(inp: std_logic_vector; old_width, delta, new_arith,
                        new_width: integer)
    return std_logic_vector
  is
    variable vec: std_logic_vector(old_width-1 downto 0);
    variable padded_inp: std_logic_vector((old_width + delta)-1  downto 0);
    variable result: std_logic_vector(new_width-1 downto 0);
  begin
    vec := inp;
    if (delta > 0) then
      padded_inp := pad_LSB(vec, old_width+delta);
      result := extend_MSB(padded_inp, new_width, new_arith);
    else
      result := extend_MSB(vec, new_width, new_arith);
    end if;
    return result;
  end;
  constant full_s_bin_pt: integer := fractional_bits(a_bin_pt, b_bin_pt);
  constant full_a_width: integer := full_s_width;
  constant full_b_width: integer := full_s_width;
  signal full_a: std_logic_vector(full_a_width - 1 downto 0);
  signal full_b: std_logic_vector(full_b_width - 1 downto 0);
  signal core_s: std_logic_vector(full_s_width - 1 downto 0);
  signal conv_s: std_logic_vector(s_width - 1 downto 0);
  signal temp_cout : std_logic;
  signal internal_clr: std_logic;
  signal internal_ce: std_logic;
  signal extra_reg_ce: std_logic;
  signal override: std_logic;
  signal logic1: std_logic_vector(0 downto 0);
  component addsb_11_0_8f54fdb6bda2d271
    port (
          a: in std_logic_vector(17 - 1 downto 0);
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(17 - 1 downto 0)
    );
  end component;
  attribute syn_black_box of addsb_11_0_8f54fdb6bda2d271:
    component is true;
  attribute fpga_dont_touch of addsb_11_0_8f54fdb6bda2d271:
    component is "true";
  attribute box_type of addsb_11_0_8f54fdb6bda2d271:
    component  is "black_box";
begin
  internal_clr <= (clr or (rst(0))) and ce;
  internal_ce <= ce and en(0);
  logic1(0) <= '1';
  addsub_process: process (a, b, core_s)
  begin
    full_a <= format_input (a, a_width, b_bin_pt - a_bin_pt, a_arith,
                            full_a_width);
    full_b <= format_input (b, b_width, a_bin_pt - b_bin_pt, b_arith,
                            full_b_width);
    conv_s <= convert_type (core_s, full_s_width, full_s_bin_pt, full_s_arith,
                            s_width, s_bin_pt, s_arith, quantization, overflow);
  end process addsub_process;

  comp0: if ((core_name0 = "addsb_11_0_8f54fdb6bda2d271")) generate
    core_instance0: addsb_11_0_8f54fdb6bda2d271
      port map (
         a => full_a,
         s => core_s,
         b => full_b
      );
  end generate;
  latency_test: if (extra_registers > 0) generate
      override_test: if (c_latency > 1) generate
       override_pipe: synth_reg
          generic map (
            width => 1,
            latency => c_latency
          )
          port map (
            i => logic1,
            ce => internal_ce,
            clr => internal_clr,
            clk => clk,
            o(0) => override);
       extra_reg_ce <= ce and en(0) and override;
      end generate override_test;
      no_override: if ((c_latency = 0) or (c_latency = 1)) generate
       extra_reg_ce <= ce and en(0);
      end generate no_override;
      extra_reg: synth_reg
        generic map (
          width => s_width,
          latency => extra_registers
        )
        port map (
          i => conv_s,
          ce => extra_reg_ce,
          clr => internal_clr,
          clk => clk,
          o => s
        );
      cout_test: if (c_has_c_out = 1) generate
      c_out_extra_reg: synth_reg
        generic map (
          width => 1,
          latency => extra_registers
        )
        port map (
          i(0) => temp_cout,
          ce => extra_reg_ce,
          clr => internal_clr,
          clk => clk,
          o => c_out
        );
      end generate cout_test;
  end generate;
  latency_s: if ((latency = 0) or (extra_registers = 0)) generate
    s <= conv_s;
  end generate latency_s;
  latency0: if (((latency = 0) or (extra_registers = 0)) and
                 (c_has_c_out = 1)) generate
    c_out(0) <= temp_cout;
  end generate latency0;
  tie_dangling_cout: if (c_has_c_out = 0) generate
    c_out <= "0";
  end generate tie_dangling_cout;
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library block_id_calc_lib;
use block_id_calc_lib.conv_pkg.all;

entity constant_0cda9054d5 is
  port (
    op : out std_logic_vector((5 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_0cda9054d5;


architecture behavior of constant_0cda9054d5 is
begin
  op <= "10010";
end behavior;


-------------------------------------------------------------------
-- System Generator version 13.2 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
library block_id_calc_lib;
use block_id_calc_lib.conv_pkg.all;
entity convert_func_call is
    generic (
        din_width    : integer := 16;
        din_bin_pt   : integer := 4;
        din_arith    : integer := xlUnsigned;
        dout_width   : integer := 8;
        dout_bin_pt  : integer := 2;
        dout_arith   : integer := xlUnsigned;
        quantization : integer := xlTruncate;
        overflow     : integer := xlWrap);
    port (
        din : in std_logic_vector (din_width-1 downto 0);
        result : out std_logic_vector (dout_width-1 downto 0));
end convert_func_call;
architecture behavior of convert_func_call is
begin
    result <= convert_type(din, din_width, din_bin_pt, din_arith,
                           dout_width, dout_bin_pt, dout_arith,
                           quantization, overflow);
end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library block_id_calc_lib;
use block_id_calc_lib.conv_pkg.all;
entity xlconvert is
    generic (
        din_width    : integer := 16;
        din_bin_pt   : integer := 4;
        din_arith    : integer := xlUnsigned;
        dout_width   : integer := 8;
        dout_bin_pt  : integer := 2;
        dout_arith   : integer := xlUnsigned;
        en_width     : integer := 1;
        en_bin_pt    : integer := 0;
        en_arith     : integer := xlUnsigned;
        bool_conversion : integer :=0;
        latency      : integer := 0;
        quantization : integer := xlTruncate;
        overflow     : integer := xlWrap);
    port (
        din : in std_logic_vector (din_width-1 downto 0);
        en  : in std_logic_vector (en_width-1 downto 0);
        ce  : in std_logic;
        clr : in std_logic;
        clk : in std_logic;
        dout : out std_logic_vector (dout_width-1 downto 0));
end xlconvert;
architecture behavior of xlconvert is
    component synth_reg
        generic (width       : integer;
                 latency     : integer);
        port (i       : in std_logic_vector(width-1 downto 0);
              ce      : in std_logic;
              clr     : in std_logic;
              clk     : in std_logic;
              o       : out std_logic_vector(width-1 downto 0));
    end component;
    component convert_func_call
        generic (
            din_width    : integer := 16;
            din_bin_pt   : integer := 4;
            din_arith    : integer := xlUnsigned;
            dout_width   : integer := 8;
            dout_bin_pt  : integer := 2;
            dout_arith   : integer := xlUnsigned;
            quantization : integer := xlTruncate;
            overflow     : integer := xlWrap);
        port (
            din : in std_logic_vector (din_width-1 downto 0);
            result : out std_logic_vector (dout_width-1 downto 0));
    end component;
    -- synopsys translate_off
    -- synopsys translate_on
    signal result : std_logic_vector(dout_width-1 downto 0);
    signal internal_ce : std_logic;
begin
    -- synopsys translate_off
    -- synopsys translate_on
    internal_ce <= ce and en(0);

    bool_conversion_generate : if (bool_conversion = 1)
    generate
      result <= din;
    end generate;
    std_conversion_generate : if (bool_conversion = 0)
    generate
      convert : convert_func_call
        generic map (
          din_width   => din_width,
          din_bin_pt  => din_bin_pt,
          din_arith   => din_arith,
          dout_width  => dout_width,
          dout_bin_pt => dout_bin_pt,
          dout_arith  => dout_arith,
          quantization => quantization,
          overflow     => overflow)
        port map (
          din => din,
          result => result);
    end generate;
    latency_test : if (latency > 0) generate
        reg : synth_reg
            generic map (
              width => dout_width,
              latency => latency
            )
            port map (
              i => result,
              ce => internal_ce,
              clr => clr,
              clk => clk,
              o => dout
            );
    end generate;
    latency0 : if (latency = 0)
    generate
        dout <= result;
    end generate latency0;
end  behavior;

-------------------------------------------------------------------
-- System Generator version 13.2 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
library block_id_calc_lib;
use block_id_calc_lib.conv_pkg.all;
entity xlcounter_free is
  generic (
    core_name0: string := "";
    op_width: integer := 5;
    op_arith: integer := xlSigned
  );
  port (
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    op: out std_logic_vector(op_width - 1 downto 0);
    up: in std_logic_vector(0 downto 0) := (others => '0');
    load: in std_logic_vector(0 downto 0) := (others => '0');
    din: in std_logic_vector(op_width - 1 downto 0) := (others => '0');
    en: in std_logic_vector(0 downto 0);
    rst: in std_logic_vector(0 downto 0)
  );
end xlcounter_free ;
architecture behavior of xlcounter_free is
  component cntr_11_0_e7514e290b172ea1
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;
  attribute syn_black_box of cntr_11_0_e7514e290b172ea1:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_e7514e290b172ea1:
    component is "true";
  attribute box_type of cntr_11_0_e7514e290b172ea1:
    component  is "black_box";
-- synopsys translate_off
  constant zeroVec: std_logic_vector(op_width - 1 downto 0) := (others => '0');
  constant oneVec: std_logic_vector(op_width - 1 downto 0) := (others => '1');
  constant zeroStr: string(1 to op_width) :=
    std_logic_vector_to_bin_string(zeroVec);
  constant oneStr: string(1 to op_width) :=
    std_logic_vector_to_bin_string(oneVec);
-- synopsys translate_on
  signal core_sinit: std_logic;
  signal core_ce: std_logic;
  signal op_net: std_logic_vector(op_width - 1 downto 0);
begin
  core_ce <= ce and en(0);
  core_sinit <= (clr or rst(0)) and ce;
  op <= op_net;
  comp0: if ((core_name0 = "cntr_11_0_e7514e290b172ea1")) generate
    core_instance0: cntr_11_0_e7514e290b172ea1
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library block_id_calc_lib;
use block_id_calc_lib.conv_pkg.all;

entity xldivider_generator_f08ad8561ebf27647140ebdb543b552e is 
  port(
    ce:in std_logic;
    clk:in std_logic;
    dividend:in std_logic_vector(15 downto 0);
    divisor:in std_logic_vector(15 downto 0);
    fractional:out std_logic_vector(15 downto 0);
    quotient:out std_logic_vector(15 downto 0);
    rfd:out std_logic
  );
end xldivider_generator_f08ad8561ebf27647140ebdb543b552e;


architecture behavior of xldivider_generator_f08ad8561ebf27647140ebdb543b552e  is
  component dv_gn_v3_0_6a34997a8a73ba6e
    port(
      ce:in std_logic;
      clk:in std_logic;
      dividend:in std_logic_vector(15 downto 0);
      divisor:in std_logic_vector(15 downto 0);
      fractional:out std_logic_vector(15 downto 0);
      quotient:out std_logic_vector(15 downto 0);
      rfd:out std_logic
    );
end component;
begin
  dv_gn_v3_0_6a34997a8a73ba6e_instance : dv_gn_v3_0_6a34997a8a73ba6e
    port map(
      ce=>ce,
      clk=>clk,
      dividend=>dividend,
      divisor=>divisor,
      fractional=>fractional,
      quotient=>quotient,
      rfd=>rfd
    );
end  behavior;


-------------------------------------------------------------------
-- System Generator version 13.2 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
library block_id_calc_lib;
use block_id_calc_lib.conv_pkg.all;
entity xlregister is
   generic (d_width          : integer := 5;
            init_value       : bit_vector := b"00");
   port (d   : in std_logic_vector (d_width-1 downto 0);
         rst : in std_logic_vector(0 downto 0) := "0";
         en  : in std_logic_vector(0 downto 0) := "1";
         ce  : in std_logic;
         clk : in std_logic;
         q   : out std_logic_vector (d_width-1 downto 0));
end xlregister;
architecture behavior of xlregister is
   component synth_reg_w_init
      generic (width      : integer;
               init_index : integer;
               init_value : bit_vector;
               latency    : integer);
      port (i   : in std_logic_vector(width-1 downto 0);
            ce  : in std_logic;
            clr : in std_logic;
            clk : in std_logic;
            o   : out std_logic_vector(width-1 downto 0));
   end component;
   -- synopsys translate_off
   signal real_d, real_q           : real;
   -- synopsys translate_on
   signal internal_clr             : std_logic;
   signal internal_ce              : std_logic;
begin
   internal_clr <= rst(0) and ce;
   internal_ce  <= en(0) and ce;
   synth_reg_inst : synth_reg_w_init
      generic map (width      => d_width,
                   init_index => 2,
                   init_value => init_value,
                   latency    => 1)
      port map (i   => d,
                ce  => internal_ce,
                clr => internal_clr,
                clk => clk,
                o   => q);
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library block_id_calc_lib;
use block_id_calc_lib.conv_pkg.all;

entity relational_02f5922aea is
  port (
    a : in std_logic_vector((8 - 1) downto 0);
    b : in std_logic_vector((5 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_02f5922aea;


architecture behavior of relational_02f5922aea is
  signal a_1_31: unsigned((8 - 1) downto 0);
  signal b_1_34: unsigned((5 - 1) downto 0);
  signal cast_12_17: unsigned((8 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_12_17 <= u2u_cast(b_1_34, 0, 8, 0);
  result_12_3_rel <= a_1_31 = cast_12_17;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
library block_id_calc_lib;
use block_id_calc_lib.conv_pkg.all;

-- Generated from Simulink block "block_id_calc"

entity block_id_calc is
  port (
    block_idx_in: in std_logic_vector(15 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    en: in std_logic; 
    grid_x_in: in std_logic_vector(15 downto 0); 
    idx_in: in std_logic_vector(15 downto 0); 
    block_id_x_out: out std_logic_vector(15 downto 0); 
    block_id_y_out: out std_logic_vector(15 downto 0); 
    valid: out std_logic
  );
end block_id_calc;

architecture structural of block_id_calc is
  attribute core_generation_info: string;
  attribute core_generation_info of structural : architecture is "block_id_calc,sysgen_core,{clock_period=10.00000000,clocking=Clock_Enables,compilation=NGC_Netlist,sample_periods=1.00000000000,testbench=1,total_blocks=28,xilinx_adder_subtracter_block=1,xilinx_arithmetic_relational_operator_block=1,xilinx_constant_block_block=1,xilinx_counter_block=1,xilinx_divider_generator_3_0_block=1,xilinx_gateway_in_block=4,xilinx_gateway_out_block=3,xilinx_register_block=4,xilinx_resource_estimator_block=1,xilinx_system_generator_block=1,xilinx_type_converter_block=1,}";

  signal addsub_s_net: std_logic_vector(15 downto 0);
  signal block_id_x_out_net: std_logic_vector(15 downto 0);
  signal block_id_y_out_net: std_logic_vector(15 downto 0);
  signal block_idx_in_net: std_logic_vector(15 downto 0);
  signal ce_1_sg_x0: std_logic;
  signal clk_1_sg_x0: std_logic;
  signal constant3_op_net: std_logic_vector(4 downto 0);
  signal convert_dout_net: std_logic;
  signal counter_op_net: std_logic_vector(7 downto 0);
  signal en_net: std_logic;
  signal grid_x_in_net: std_logic_vector(15 downto 0);
  signal idx_in_net: std_logic_vector(15 downto 0);
  signal register1_q_net: std_logic_vector(15 downto 0);
  signal register2_q_net: std_logic_vector(15 downto 0);
  signal register3_q_net: std_logic;
  signal register_q_net: std_logic_vector(15 downto 0);
  signal valid_net: std_logic;

begin
  block_idx_in_net <= block_idx_in;
  ce_1_sg_x0 <= ce_1;
  clk_1_sg_x0 <= clk_1;
  en_net <= en;
  grid_x_in_net <= grid_x_in;
  idx_in_net <= idx_in;
  block_id_x_out <= block_id_x_out_net;
  block_id_y_out <= block_id_y_out_net;
  valid <= valid_net;

  addsub: entity block_id_calc_lib.xladdsub
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 16,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 16,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 17,
      core_name0 => "addsb_11_0_8f54fdb6bda2d271",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 17,
      latency => 0,
      overflow => 2,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 16
    )
    port map (
      a => register_q_net,
      b => register1_q_net,
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      en => "1",
      s => addsub_s_net
    );

  constant3: entity block_id_calc_lib.constant_0cda9054d5
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant3_op_net
    );

  convert: entity block_id_calc_lib.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      din(0) => en_net,
      en => "1",
      dout(0) => convert_dout_net
    );

  counter: entity block_id_calc_lib.xlcounter_free
    generic map (
      core_name0 => "cntr_11_0_e7514e290b172ea1",
      op_arith => xlUnsigned,
      op_width => 8
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      en(0) => register3_q_net,
      rst(0) => valid_net,
      op => counter_op_net
    );

  divider_generator_3_0: entity block_id_calc_lib.xldivider_generator_f08ad8561ebf27647140ebdb543b552e
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      dividend => addsub_s_net,
      divisor => register2_q_net,
      fractional => block_id_x_out_net,
      quotient => block_id_y_out_net
    );

  register1: entity block_id_calc_lib.xlregister
    generic map (
      d_width => 16,
      init_value => b"0000000000000000"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d => idx_in_net,
      en(0) => convert_dout_net,
      rst => "0",
      q => register1_q_net
    );

  register2: entity block_id_calc_lib.xlregister
    generic map (
      d_width => 16,
      init_value => b"0000000000000000"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d => grid_x_in_net,
      en(0) => convert_dout_net,
      rst => "0",
      q => register2_q_net
    );

  register3: entity block_id_calc_lib.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d(0) => convert_dout_net,
      en(0) => convert_dout_net,
      rst(0) => valid_net,
      q(0) => register3_q_net
    );

  register_x0: entity block_id_calc_lib.xlregister
    generic map (
      d_width => 16,
      init_value => b"0000000000000000"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d => block_idx_in_net,
      en(0) => convert_dout_net,
      rst => "0",
      q => register_q_net
    );

  relational: entity block_id_calc_lib.relational_02f5922aea
    port map (
      a => counter_op_net,
      b => constant3_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => valid_net
    );

end structural;
