--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2012 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_84fc5d4200208b4e.vhd when simulating
-- the core, addsb_11_0_84fc5d4200208b4e. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_84fc5d4200208b4e IS
  PORT (
    a : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
  );
END addsb_11_0_84fc5d4200208b4e;

ARCHITECTURE addsb_11_0_84fc5d4200208b4e_a OF addsb_11_0_84fc5d4200208b4e IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_84fc5d4200208b4e
  PORT (
    a : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_84fc5d4200208b4e USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 1,
      c_a_width => 7,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 1,
      c_b_value => "0000000",
      c_b_width => 7,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 0,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 0,
      c_out_width => 7,
      c_sclr_overrides_sset => 0,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_84fc5d4200208b4e
  PORT MAP (
    a => a,
    b => b,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_84fc5d4200208b4e_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2012 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_e7514e290b172ea1.vhd when simulating
-- the core, cntr_11_0_e7514e290b172ea1. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_e7514e290b172ea1 IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END cntr_11_0_e7514e290b172ea1;

ARCHITECTURE cntr_11_0_e7514e290b172ea1_a OF cntr_11_0_e7514e290b172ea1 IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_e7514e290b172ea1
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_e7514e290b172ea1 USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 8,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_e7514e290b172ea1
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_e7514e290b172ea1_a;
--------------------------------------------------------------------------------
-- Copyright (c) 1995-2011 Xilinx, Inc.  All rights reserved.
--------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version: O.61xd
--  \   \         Application: netgen
--  /   /         Filename: dv_gn_v3_0_c648497ecac7f882.vhd
-- /___/   /\     Timestamp: Thu Apr 12 11:30:55 2012
-- \   \  /  \ 
--  \___\/\___\
--             
-- Command	: -intstyle ise -w -sim -ofmt vhdl ./tmp/_cg/dv_gn_v3_0_c648497ecac7f882.ngc ./tmp/_cg/dv_gn_v3_0_c648497ecac7f882.vhd 
-- Device	: 6vcx75tff484-2
-- Input file	: ./tmp/_cg/dv_gn_v3_0_c648497ecac7f882.ngc
-- Output file	: ./tmp/_cg/dv_gn_v3_0_c648497ecac7f882.vhd
-- # of Entities	: 1
-- Design Name	: dv_gn_v3_0_c648497ecac7f882
-- Xilinx	: c:\xilinx\13.2\ise_ds\ise\
--             
-- Purpose:    
--     This VHDL netlist is a verification model and uses simulation 
--     primitives which may not represent the true implementation of the 
--     device, however the netlist is functionally correct and should not 
--     be modified. This file cannot be synthesized and should only be used 
--     with supported simulation tools.
--             
-- Reference:  
--     Command Line Tools User Guide, Chapter 23
--     Synthesis and Simulation Design Guide, Chapter 6
--             
--------------------------------------------------------------------------------


-- synthesis translate_off
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;
use UNISIM.VPKG.ALL;

entity dv_gn_v3_0_c648497ecac7f882 is
  port (
    ce : in STD_LOGIC := 'X'; 
    rfd : out STD_LOGIC; 
    clk : in STD_LOGIC := 'X'; 
    dividend : in STD_LOGIC_VECTOR ( 11 downto 0 ); 
    quotient : out STD_LOGIC_VECTOR ( 11 downto 0 ); 
    divisor : in STD_LOGIC_VECTOR ( 5 downto 0 ); 
    fractional : out STD_LOGIC_VECTOR ( 15 downto 0 ) 
  );
end dv_gn_v3_0_c648497ecac7f882;

architecture STRUCTURE of dv_gn_v3_0_c648497ecac7f882 is
  signal NlwRenamedSig_OI_rfd : STD_LOGIC; 
  signal blk00000003_sig000005e5 : STD_LOGIC; 
  signal blk00000003_sig000005e4 : STD_LOGIC; 
  signal blk00000003_sig000005e3 : STD_LOGIC; 
  signal blk00000003_sig000005e2 : STD_LOGIC; 
  signal blk00000003_sig000005e1 : STD_LOGIC; 
  signal blk00000003_sig000005e0 : STD_LOGIC; 
  signal blk00000003_sig000005df : STD_LOGIC; 
  signal blk00000003_sig000005de : STD_LOGIC; 
  signal blk00000003_sig000005dd : STD_LOGIC; 
  signal blk00000003_sig000005dc : STD_LOGIC; 
  signal blk00000003_sig000005db : STD_LOGIC; 
  signal blk00000003_sig000005da : STD_LOGIC; 
  signal blk00000003_sig000005d9 : STD_LOGIC; 
  signal blk00000003_sig000005d8 : STD_LOGIC; 
  signal blk00000003_sig000005d7 : STD_LOGIC; 
  signal blk00000003_sig000005d6 : STD_LOGIC; 
  signal blk00000003_sig000005d5 : STD_LOGIC; 
  signal blk00000003_sig000005d4 : STD_LOGIC; 
  signal blk00000003_sig000005d3 : STD_LOGIC; 
  signal blk00000003_sig000005d2 : STD_LOGIC; 
  signal blk00000003_sig000005d1 : STD_LOGIC; 
  signal blk00000003_sig000005d0 : STD_LOGIC; 
  signal blk00000003_sig000005cf : STD_LOGIC; 
  signal blk00000003_sig000005ce : STD_LOGIC; 
  signal blk00000003_sig000005cd : STD_LOGIC; 
  signal blk00000003_sig000005cc : STD_LOGIC; 
  signal blk00000003_sig000005cb : STD_LOGIC; 
  signal blk00000003_sig000005ca : STD_LOGIC; 
  signal blk00000003_sig000005c9 : STD_LOGIC; 
  signal blk00000003_sig000005c8 : STD_LOGIC; 
  signal blk00000003_sig000005c7 : STD_LOGIC; 
  signal blk00000003_sig000005c6 : STD_LOGIC; 
  signal blk00000003_sig000005c5 : STD_LOGIC; 
  signal blk00000003_sig000005c4 : STD_LOGIC; 
  signal blk00000003_sig000005c3 : STD_LOGIC; 
  signal blk00000003_sig000005c2 : STD_LOGIC; 
  signal blk00000003_sig000005c1 : STD_LOGIC; 
  signal blk00000003_sig000005c0 : STD_LOGIC; 
  signal blk00000003_sig000005bf : STD_LOGIC; 
  signal blk00000003_sig000005be : STD_LOGIC; 
  signal blk00000003_sig000005bd : STD_LOGIC; 
  signal blk00000003_sig000005bc : STD_LOGIC; 
  signal blk00000003_sig000005bb : STD_LOGIC; 
  signal blk00000003_sig000005ba : STD_LOGIC; 
  signal blk00000003_sig000005b9 : STD_LOGIC; 
  signal blk00000003_sig000005b8 : STD_LOGIC; 
  signal blk00000003_sig000005b7 : STD_LOGIC; 
  signal blk00000003_sig000005b6 : STD_LOGIC; 
  signal blk00000003_sig000005b5 : STD_LOGIC; 
  signal blk00000003_sig000005b4 : STD_LOGIC; 
  signal blk00000003_sig000005b3 : STD_LOGIC; 
  signal blk00000003_sig000005b2 : STD_LOGIC; 
  signal blk00000003_sig000005b1 : STD_LOGIC; 
  signal blk00000003_sig000005b0 : STD_LOGIC; 
  signal blk00000003_sig000005af : STD_LOGIC; 
  signal blk00000003_sig000005ae : STD_LOGIC; 
  signal blk00000003_sig000005ad : STD_LOGIC; 
  signal blk00000003_sig000005ac : STD_LOGIC; 
  signal blk00000003_sig000005ab : STD_LOGIC; 
  signal blk00000003_sig000005aa : STD_LOGIC; 
  signal blk00000003_sig000005a9 : STD_LOGIC; 
  signal blk00000003_sig000005a8 : STD_LOGIC; 
  signal blk00000003_sig000005a7 : STD_LOGIC; 
  signal blk00000003_sig000005a6 : STD_LOGIC; 
  signal blk00000003_sig000005a5 : STD_LOGIC; 
  signal blk00000003_sig000005a4 : STD_LOGIC; 
  signal blk00000003_sig000005a3 : STD_LOGIC; 
  signal blk00000003_sig000005a2 : STD_LOGIC; 
  signal blk00000003_sig000005a1 : STD_LOGIC; 
  signal blk00000003_sig000005a0 : STD_LOGIC; 
  signal blk00000003_sig0000059f : STD_LOGIC; 
  signal blk00000003_sig0000059e : STD_LOGIC; 
  signal blk00000003_sig0000059d : STD_LOGIC; 
  signal blk00000003_sig0000059c : STD_LOGIC; 
  signal blk00000003_sig0000059b : STD_LOGIC; 
  signal blk00000003_sig0000059a : STD_LOGIC; 
  signal blk00000003_sig00000599 : STD_LOGIC; 
  signal blk00000003_sig00000598 : STD_LOGIC; 
  signal blk00000003_sig00000597 : STD_LOGIC; 
  signal blk00000003_sig00000596 : STD_LOGIC; 
  signal blk00000003_sig00000595 : STD_LOGIC; 
  signal blk00000003_sig00000594 : STD_LOGIC; 
  signal blk00000003_sig00000593 : STD_LOGIC; 
  signal blk00000003_sig00000592 : STD_LOGIC; 
  signal blk00000003_sig00000591 : STD_LOGIC; 
  signal blk00000003_sig00000590 : STD_LOGIC; 
  signal blk00000003_sig0000058f : STD_LOGIC; 
  signal blk00000003_sig0000058e : STD_LOGIC; 
  signal blk00000003_sig0000058d : STD_LOGIC; 
  signal blk00000003_sig0000058c : STD_LOGIC; 
  signal blk00000003_sig0000058b : STD_LOGIC; 
  signal blk00000003_sig0000058a : STD_LOGIC; 
  signal blk00000003_sig00000589 : STD_LOGIC; 
  signal blk00000003_sig00000588 : STD_LOGIC; 
  signal blk00000003_sig00000587 : STD_LOGIC; 
  signal blk00000003_sig00000586 : STD_LOGIC; 
  signal blk00000003_sig00000585 : STD_LOGIC; 
  signal blk00000003_sig00000584 : STD_LOGIC; 
  signal blk00000003_sig00000583 : STD_LOGIC; 
  signal blk00000003_sig00000582 : STD_LOGIC; 
  signal blk00000003_sig00000581 : STD_LOGIC; 
  signal blk00000003_sig00000580 : STD_LOGIC; 
  signal blk00000003_sig0000057f : STD_LOGIC; 
  signal blk00000003_sig0000057e : STD_LOGIC; 
  signal blk00000003_sig0000057d : STD_LOGIC; 
  signal blk00000003_sig0000057c : STD_LOGIC; 
  signal blk00000003_sig0000057b : STD_LOGIC; 
  signal blk00000003_sig0000057a : STD_LOGIC; 
  signal blk00000003_sig00000579 : STD_LOGIC; 
  signal blk00000003_sig00000578 : STD_LOGIC; 
  signal blk00000003_sig00000577 : STD_LOGIC; 
  signal blk00000003_sig00000576 : STD_LOGIC; 
  signal blk00000003_sig00000575 : STD_LOGIC; 
  signal blk00000003_sig00000574 : STD_LOGIC; 
  signal blk00000003_sig00000573 : STD_LOGIC; 
  signal blk00000003_sig00000572 : STD_LOGIC; 
  signal blk00000003_sig00000571 : STD_LOGIC; 
  signal blk00000003_sig00000570 : STD_LOGIC; 
  signal blk00000003_sig0000056f : STD_LOGIC; 
  signal blk00000003_sig0000056e : STD_LOGIC; 
  signal blk00000003_sig0000056d : STD_LOGIC; 
  signal blk00000003_sig0000056c : STD_LOGIC; 
  signal blk00000003_sig0000056b : STD_LOGIC; 
  signal blk00000003_sig0000056a : STD_LOGIC; 
  signal blk00000003_sig00000569 : STD_LOGIC; 
  signal blk00000003_sig00000568 : STD_LOGIC; 
  signal blk00000003_sig00000567 : STD_LOGIC; 
  signal blk00000003_sig00000566 : STD_LOGIC; 
  signal blk00000003_sig00000565 : STD_LOGIC; 
  signal blk00000003_sig00000564 : STD_LOGIC; 
  signal blk00000003_sig00000563 : STD_LOGIC; 
  signal blk00000003_sig00000562 : STD_LOGIC; 
  signal blk00000003_sig00000561 : STD_LOGIC; 
  signal blk00000003_sig00000560 : STD_LOGIC; 
  signal blk00000003_sig0000055f : STD_LOGIC; 
  signal blk00000003_sig0000055e : STD_LOGIC; 
  signal blk00000003_sig0000055d : STD_LOGIC; 
  signal blk00000003_sig0000055c : STD_LOGIC; 
  signal blk00000003_sig0000055b : STD_LOGIC; 
  signal blk00000003_sig0000055a : STD_LOGIC; 
  signal blk00000003_sig00000559 : STD_LOGIC; 
  signal blk00000003_sig00000558 : STD_LOGIC; 
  signal blk00000003_sig00000557 : STD_LOGIC; 
  signal blk00000003_sig00000556 : STD_LOGIC; 
  signal blk00000003_sig00000555 : STD_LOGIC; 
  signal blk00000003_sig00000554 : STD_LOGIC; 
  signal blk00000003_sig00000553 : STD_LOGIC; 
  signal blk00000003_sig00000552 : STD_LOGIC; 
  signal blk00000003_sig00000551 : STD_LOGIC; 
  signal blk00000003_sig00000550 : STD_LOGIC; 
  signal blk00000003_sig0000054f : STD_LOGIC; 
  signal blk00000003_sig0000054e : STD_LOGIC; 
  signal blk00000003_sig0000054d : STD_LOGIC; 
  signal blk00000003_sig0000054c : STD_LOGIC; 
  signal blk00000003_sig0000054b : STD_LOGIC; 
  signal blk00000003_sig0000054a : STD_LOGIC; 
  signal blk00000003_sig00000549 : STD_LOGIC; 
  signal blk00000003_sig00000548 : STD_LOGIC; 
  signal blk00000003_sig00000547 : STD_LOGIC; 
  signal blk00000003_sig00000546 : STD_LOGIC; 
  signal blk00000003_sig00000545 : STD_LOGIC; 
  signal blk00000003_sig00000544 : STD_LOGIC; 
  signal blk00000003_sig00000543 : STD_LOGIC; 
  signal blk00000003_sig00000542 : STD_LOGIC; 
  signal blk00000003_sig00000541 : STD_LOGIC; 
  signal blk00000003_sig00000540 : STD_LOGIC; 
  signal blk00000003_sig0000053f : STD_LOGIC; 
  signal blk00000003_sig0000053e : STD_LOGIC; 
  signal blk00000003_sig0000053d : STD_LOGIC; 
  signal blk00000003_sig0000053c : STD_LOGIC; 
  signal blk00000003_sig0000053b : STD_LOGIC; 
  signal blk00000003_sig0000053a : STD_LOGIC; 
  signal blk00000003_sig00000539 : STD_LOGIC; 
  signal blk00000003_sig00000538 : STD_LOGIC; 
  signal blk00000003_sig00000537 : STD_LOGIC; 
  signal blk00000003_sig00000536 : STD_LOGIC; 
  signal blk00000003_sig00000535 : STD_LOGIC; 
  signal blk00000003_sig00000534 : STD_LOGIC; 
  signal blk00000003_sig00000533 : STD_LOGIC; 
  signal blk00000003_sig00000532 : STD_LOGIC; 
  signal blk00000003_sig00000531 : STD_LOGIC; 
  signal blk00000003_sig00000530 : STD_LOGIC; 
  signal blk00000003_sig0000052f : STD_LOGIC; 
  signal blk00000003_sig0000052e : STD_LOGIC; 
  signal blk00000003_sig0000052d : STD_LOGIC; 
  signal blk00000003_sig0000052c : STD_LOGIC; 
  signal blk00000003_sig0000052b : STD_LOGIC; 
  signal blk00000003_sig0000052a : STD_LOGIC; 
  signal blk00000003_sig00000529 : STD_LOGIC; 
  signal blk00000003_sig00000528 : STD_LOGIC; 
  signal blk00000003_sig00000527 : STD_LOGIC; 
  signal blk00000003_sig00000526 : STD_LOGIC; 
  signal blk00000003_sig00000525 : STD_LOGIC; 
  signal blk00000003_sig00000524 : STD_LOGIC; 
  signal blk00000003_sig00000523 : STD_LOGIC; 
  signal blk00000003_sig00000522 : STD_LOGIC; 
  signal blk00000003_sig00000521 : STD_LOGIC; 
  signal blk00000003_sig00000520 : STD_LOGIC; 
  signal blk00000003_sig0000051f : STD_LOGIC; 
  signal blk00000003_sig0000051e : STD_LOGIC; 
  signal blk00000003_sig0000051d : STD_LOGIC; 
  signal blk00000003_sig0000051c : STD_LOGIC; 
  signal blk00000003_sig0000051b : STD_LOGIC; 
  signal blk00000003_sig0000051a : STD_LOGIC; 
  signal blk00000003_sig00000519 : STD_LOGIC; 
  signal blk00000003_sig00000518 : STD_LOGIC; 
  signal blk00000003_sig00000517 : STD_LOGIC; 
  signal blk00000003_sig00000516 : STD_LOGIC; 
  signal blk00000003_sig00000515 : STD_LOGIC; 
  signal blk00000003_sig00000514 : STD_LOGIC; 
  signal blk00000003_sig00000513 : STD_LOGIC; 
  signal blk00000003_sig00000512 : STD_LOGIC; 
  signal blk00000003_sig00000511 : STD_LOGIC; 
  signal blk00000003_sig00000510 : STD_LOGIC; 
  signal blk00000003_sig0000050f : STD_LOGIC; 
  signal blk00000003_sig0000050e : STD_LOGIC; 
  signal blk00000003_sig0000050d : STD_LOGIC; 
  signal blk00000003_sig0000050c : STD_LOGIC; 
  signal blk00000003_sig0000050b : STD_LOGIC; 
  signal blk00000003_sig0000050a : STD_LOGIC; 
  signal blk00000003_sig00000509 : STD_LOGIC; 
  signal blk00000003_sig00000508 : STD_LOGIC; 
  signal blk00000003_sig00000507 : STD_LOGIC; 
  signal blk00000003_sig00000506 : STD_LOGIC; 
  signal blk00000003_sig00000505 : STD_LOGIC; 
  signal blk00000003_sig00000504 : STD_LOGIC; 
  signal blk00000003_sig00000503 : STD_LOGIC; 
  signal blk00000003_sig00000502 : STD_LOGIC; 
  signal blk00000003_sig00000501 : STD_LOGIC; 
  signal blk00000003_sig00000500 : STD_LOGIC; 
  signal blk00000003_sig000004ff : STD_LOGIC; 
  signal blk00000003_sig000004fe : STD_LOGIC; 
  signal blk00000003_sig000004fd : STD_LOGIC; 
  signal blk00000003_sig000004fc : STD_LOGIC; 
  signal blk00000003_sig000004fb : STD_LOGIC; 
  signal blk00000003_sig000004fa : STD_LOGIC; 
  signal blk00000003_sig000004f9 : STD_LOGIC; 
  signal blk00000003_sig000004f8 : STD_LOGIC; 
  signal blk00000003_sig000004f7 : STD_LOGIC; 
  signal blk00000003_sig000004f6 : STD_LOGIC; 
  signal blk00000003_sig000004f5 : STD_LOGIC; 
  signal blk00000003_sig000004f4 : STD_LOGIC; 
  signal blk00000003_sig000004f3 : STD_LOGIC; 
  signal blk00000003_sig000004f2 : STD_LOGIC; 
  signal blk00000003_sig000004f1 : STD_LOGIC; 
  signal blk00000003_sig000004f0 : STD_LOGIC; 
  signal blk00000003_sig000004ef : STD_LOGIC; 
  signal blk00000003_sig000004ee : STD_LOGIC; 
  signal blk00000003_sig000004ed : STD_LOGIC; 
  signal blk00000003_sig000004ec : STD_LOGIC; 
  signal blk00000003_sig000004eb : STD_LOGIC; 
  signal blk00000003_sig000004ea : STD_LOGIC; 
  signal blk00000003_sig000004e9 : STD_LOGIC; 
  signal blk00000003_sig000004e8 : STD_LOGIC; 
  signal blk00000003_sig000004e7 : STD_LOGIC; 
  signal blk00000003_sig000004e6 : STD_LOGIC; 
  signal blk00000003_sig000004e5 : STD_LOGIC; 
  signal blk00000003_sig000004e4 : STD_LOGIC; 
  signal blk00000003_sig000004e3 : STD_LOGIC; 
  signal blk00000003_sig000004e2 : STD_LOGIC; 
  signal blk00000003_sig000004e1 : STD_LOGIC; 
  signal blk00000003_sig000004e0 : STD_LOGIC; 
  signal blk00000003_sig000004df : STD_LOGIC; 
  signal blk00000003_sig000004de : STD_LOGIC; 
  signal blk00000003_sig000004dd : STD_LOGIC; 
  signal blk00000003_sig000004dc : STD_LOGIC; 
  signal blk00000003_sig000004db : STD_LOGIC; 
  signal blk00000003_sig000004da : STD_LOGIC; 
  signal blk00000003_sig000004d9 : STD_LOGIC; 
  signal blk00000003_sig000004d8 : STD_LOGIC; 
  signal blk00000003_sig000004d7 : STD_LOGIC; 
  signal blk00000003_sig000004d6 : STD_LOGIC; 
  signal blk00000003_sig000004d5 : STD_LOGIC; 
  signal blk00000003_sig000004d4 : STD_LOGIC; 
  signal blk00000003_sig000004d3 : STD_LOGIC; 
  signal blk00000003_sig000004d2 : STD_LOGIC; 
  signal blk00000003_sig000004d1 : STD_LOGIC; 
  signal blk00000003_sig000004d0 : STD_LOGIC; 
  signal blk00000003_sig000004cf : STD_LOGIC; 
  signal blk00000003_sig000004ce : STD_LOGIC; 
  signal blk00000003_sig000004cd : STD_LOGIC; 
  signal blk00000003_sig000004cc : STD_LOGIC; 
  signal blk00000003_sig000004cb : STD_LOGIC; 
  signal blk00000003_sig000004ca : STD_LOGIC; 
  signal blk00000003_sig000004c9 : STD_LOGIC; 
  signal blk00000003_sig000004c8 : STD_LOGIC; 
  signal blk00000003_sig000004c7 : STD_LOGIC; 
  signal blk00000003_sig000004c6 : STD_LOGIC; 
  signal blk00000003_sig000004c5 : STD_LOGIC; 
  signal blk00000003_sig000004c4 : STD_LOGIC; 
  signal blk00000003_sig000004c3 : STD_LOGIC; 
  signal blk00000003_sig000004c2 : STD_LOGIC; 
  signal blk00000003_sig000004c1 : STD_LOGIC; 
  signal blk00000003_sig000004c0 : STD_LOGIC; 
  signal blk00000003_sig000004bf : STD_LOGIC; 
  signal blk00000003_sig000004be : STD_LOGIC; 
  signal blk00000003_sig000004bd : STD_LOGIC; 
  signal blk00000003_sig000004bc : STD_LOGIC; 
  signal blk00000003_sig000004bb : STD_LOGIC; 
  signal blk00000003_sig000004ba : STD_LOGIC; 
  signal blk00000003_sig000004b9 : STD_LOGIC; 
  signal blk00000003_sig000004b8 : STD_LOGIC; 
  signal blk00000003_sig000004b7 : STD_LOGIC; 
  signal blk00000003_sig000004b6 : STD_LOGIC; 
  signal blk00000003_sig000004b5 : STD_LOGIC; 
  signal blk00000003_sig000004b4 : STD_LOGIC; 
  signal blk00000003_sig000004b3 : STD_LOGIC; 
  signal blk00000003_sig000004b2 : STD_LOGIC; 
  signal blk00000003_sig000004b1 : STD_LOGIC; 
  signal blk00000003_sig000004b0 : STD_LOGIC; 
  signal blk00000003_sig000004af : STD_LOGIC; 
  signal blk00000003_sig000004ae : STD_LOGIC; 
  signal blk00000003_sig000004ad : STD_LOGIC; 
  signal blk00000003_sig000004ac : STD_LOGIC; 
  signal blk00000003_sig000004ab : STD_LOGIC; 
  signal blk00000003_sig000004aa : STD_LOGIC; 
  signal blk00000003_sig000004a9 : STD_LOGIC; 
  signal blk00000003_sig000004a8 : STD_LOGIC; 
  signal blk00000003_sig000004a7 : STD_LOGIC; 
  signal blk00000003_sig000004a6 : STD_LOGIC; 
  signal blk00000003_sig000004a5 : STD_LOGIC; 
  signal blk00000003_sig000004a4 : STD_LOGIC; 
  signal blk00000003_sig000004a3 : STD_LOGIC; 
  signal blk00000003_sig000004a2 : STD_LOGIC; 
  signal blk00000003_sig000004a1 : STD_LOGIC; 
  signal blk00000003_sig000004a0 : STD_LOGIC; 
  signal blk00000003_sig0000049f : STD_LOGIC; 
  signal blk00000003_sig0000049e : STD_LOGIC; 
  signal blk00000003_sig0000049d : STD_LOGIC; 
  signal blk00000003_sig0000049c : STD_LOGIC; 
  signal blk00000003_sig0000049b : STD_LOGIC; 
  signal blk00000003_sig0000049a : STD_LOGIC; 
  signal blk00000003_sig00000499 : STD_LOGIC; 
  signal blk00000003_sig00000498 : STD_LOGIC; 
  signal blk00000003_sig00000497 : STD_LOGIC; 
  signal blk00000003_sig00000496 : STD_LOGIC; 
  signal blk00000003_sig00000495 : STD_LOGIC; 
  signal blk00000003_sig00000494 : STD_LOGIC; 
  signal blk00000003_sig00000493 : STD_LOGIC; 
  signal blk00000003_sig00000492 : STD_LOGIC; 
  signal blk00000003_sig00000491 : STD_LOGIC; 
  signal blk00000003_sig00000490 : STD_LOGIC; 
  signal blk00000003_sig0000048f : STD_LOGIC; 
  signal blk00000003_sig0000048e : STD_LOGIC; 
  signal blk00000003_sig0000048d : STD_LOGIC; 
  signal blk00000003_sig0000048c : STD_LOGIC; 
  signal blk00000003_sig0000048b : STD_LOGIC; 
  signal blk00000003_sig0000048a : STD_LOGIC; 
  signal blk00000003_sig00000489 : STD_LOGIC; 
  signal blk00000003_sig00000488 : STD_LOGIC; 
  signal blk00000003_sig00000487 : STD_LOGIC; 
  signal blk00000003_sig00000486 : STD_LOGIC; 
  signal blk00000003_sig00000485 : STD_LOGIC; 
  signal blk00000003_sig00000484 : STD_LOGIC; 
  signal blk00000003_sig00000483 : STD_LOGIC; 
  signal blk00000003_sig00000482 : STD_LOGIC; 
  signal blk00000003_sig00000481 : STD_LOGIC; 
  signal blk00000003_sig00000480 : STD_LOGIC; 
  signal blk00000003_sig0000047f : STD_LOGIC; 
  signal blk00000003_sig0000047e : STD_LOGIC; 
  signal blk00000003_sig0000047d : STD_LOGIC; 
  signal blk00000003_sig0000047c : STD_LOGIC; 
  signal blk00000003_sig0000047b : STD_LOGIC; 
  signal blk00000003_sig0000047a : STD_LOGIC; 
  signal blk00000003_sig00000479 : STD_LOGIC; 
  signal blk00000003_sig00000478 : STD_LOGIC; 
  signal blk00000003_sig00000477 : STD_LOGIC; 
  signal blk00000003_sig00000476 : STD_LOGIC; 
  signal blk00000003_sig00000475 : STD_LOGIC; 
  signal blk00000003_sig00000474 : STD_LOGIC; 
  signal blk00000003_sig00000473 : STD_LOGIC; 
  signal blk00000003_sig00000472 : STD_LOGIC; 
  signal blk00000003_sig00000471 : STD_LOGIC; 
  signal blk00000003_sig00000470 : STD_LOGIC; 
  signal blk00000003_sig0000046f : STD_LOGIC; 
  signal blk00000003_sig0000046e : STD_LOGIC; 
  signal blk00000003_sig0000046d : STD_LOGIC; 
  signal blk00000003_sig0000046c : STD_LOGIC; 
  signal blk00000003_sig0000046b : STD_LOGIC; 
  signal blk00000003_sig0000046a : STD_LOGIC; 
  signal blk00000003_sig00000469 : STD_LOGIC; 
  signal blk00000003_sig00000468 : STD_LOGIC; 
  signal blk00000003_sig00000467 : STD_LOGIC; 
  signal blk00000003_sig00000466 : STD_LOGIC; 
  signal blk00000003_sig00000465 : STD_LOGIC; 
  signal blk00000003_sig00000464 : STD_LOGIC; 
  signal blk00000003_sig00000463 : STD_LOGIC; 
  signal blk00000003_sig00000462 : STD_LOGIC; 
  signal blk00000003_sig00000461 : STD_LOGIC; 
  signal blk00000003_sig00000460 : STD_LOGIC; 
  signal blk00000003_sig0000045f : STD_LOGIC; 
  signal blk00000003_sig0000045e : STD_LOGIC; 
  signal blk00000003_sig0000045d : STD_LOGIC; 
  signal blk00000003_sig0000045c : STD_LOGIC; 
  signal blk00000003_sig0000045b : STD_LOGIC; 
  signal blk00000003_sig0000045a : STD_LOGIC; 
  signal blk00000003_sig00000459 : STD_LOGIC; 
  signal blk00000003_sig00000458 : STD_LOGIC; 
  signal blk00000003_sig00000457 : STD_LOGIC; 
  signal blk00000003_sig00000456 : STD_LOGIC; 
  signal blk00000003_sig00000455 : STD_LOGIC; 
  signal blk00000003_sig00000454 : STD_LOGIC; 
  signal blk00000003_sig00000453 : STD_LOGIC; 
  signal blk00000003_sig00000452 : STD_LOGIC; 
  signal blk00000003_sig00000451 : STD_LOGIC; 
  signal blk00000003_sig00000450 : STD_LOGIC; 
  signal blk00000003_sig0000044f : STD_LOGIC; 
  signal blk00000003_sig0000044e : STD_LOGIC; 
  signal blk00000003_sig0000044d : STD_LOGIC; 
  signal blk00000003_sig0000044c : STD_LOGIC; 
  signal blk00000003_sig0000044b : STD_LOGIC; 
  signal blk00000003_sig0000044a : STD_LOGIC; 
  signal blk00000003_sig00000449 : STD_LOGIC; 
  signal blk00000003_sig00000448 : STD_LOGIC; 
  signal blk00000003_sig00000447 : STD_LOGIC; 
  signal blk00000003_sig00000446 : STD_LOGIC; 
  signal blk00000003_sig00000445 : STD_LOGIC; 
  signal blk00000003_sig00000444 : STD_LOGIC; 
  signal blk00000003_sig00000443 : STD_LOGIC; 
  signal blk00000003_sig00000442 : STD_LOGIC; 
  signal blk00000003_sig00000441 : STD_LOGIC; 
  signal blk00000003_sig00000440 : STD_LOGIC; 
  signal blk00000003_sig0000043f : STD_LOGIC; 
  signal blk00000003_sig0000043e : STD_LOGIC; 
  signal blk00000003_sig0000043d : STD_LOGIC; 
  signal blk00000003_sig0000043c : STD_LOGIC; 
  signal blk00000003_sig0000043b : STD_LOGIC; 
  signal blk00000003_sig0000043a : STD_LOGIC; 
  signal blk00000003_sig00000439 : STD_LOGIC; 
  signal blk00000003_sig00000438 : STD_LOGIC; 
  signal blk00000003_sig00000437 : STD_LOGIC; 
  signal blk00000003_sig00000436 : STD_LOGIC; 
  signal blk00000003_sig00000435 : STD_LOGIC; 
  signal blk00000003_sig00000434 : STD_LOGIC; 
  signal blk00000003_sig00000433 : STD_LOGIC; 
  signal blk00000003_sig00000432 : STD_LOGIC; 
  signal blk00000003_sig00000431 : STD_LOGIC; 
  signal blk00000003_sig00000430 : STD_LOGIC; 
  signal blk00000003_sig0000042f : STD_LOGIC; 
  signal blk00000003_sig0000042e : STD_LOGIC; 
  signal blk00000003_sig0000042d : STD_LOGIC; 
  signal blk00000003_sig0000042c : STD_LOGIC; 
  signal blk00000003_sig0000042b : STD_LOGIC; 
  signal blk00000003_sig0000042a : STD_LOGIC; 
  signal blk00000003_sig00000429 : STD_LOGIC; 
  signal blk00000003_sig00000428 : STD_LOGIC; 
  signal blk00000003_sig00000427 : STD_LOGIC; 
  signal blk00000003_sig00000426 : STD_LOGIC; 
  signal blk00000003_sig00000425 : STD_LOGIC; 
  signal blk00000003_sig00000424 : STD_LOGIC; 
  signal blk00000003_sig00000423 : STD_LOGIC; 
  signal blk00000003_sig00000422 : STD_LOGIC; 
  signal blk00000003_sig00000421 : STD_LOGIC; 
  signal blk00000003_sig00000420 : STD_LOGIC; 
  signal blk00000003_sig0000041f : STD_LOGIC; 
  signal blk00000003_sig0000041e : STD_LOGIC; 
  signal blk00000003_sig0000041d : STD_LOGIC; 
  signal blk00000003_sig0000041c : STD_LOGIC; 
  signal blk00000003_sig0000041b : STD_LOGIC; 
  signal blk00000003_sig0000041a : STD_LOGIC; 
  signal blk00000003_sig00000419 : STD_LOGIC; 
  signal blk00000003_sig00000418 : STD_LOGIC; 
  signal blk00000003_sig00000417 : STD_LOGIC; 
  signal blk00000003_sig00000416 : STD_LOGIC; 
  signal blk00000003_sig00000415 : STD_LOGIC; 
  signal blk00000003_sig00000414 : STD_LOGIC; 
  signal blk00000003_sig00000413 : STD_LOGIC; 
  signal blk00000003_sig00000412 : STD_LOGIC; 
  signal blk00000003_sig00000411 : STD_LOGIC; 
  signal blk00000003_sig00000410 : STD_LOGIC; 
  signal blk00000003_sig0000040f : STD_LOGIC; 
  signal blk00000003_sig0000040e : STD_LOGIC; 
  signal blk00000003_sig0000040d : STD_LOGIC; 
  signal blk00000003_sig0000040c : STD_LOGIC; 
  signal blk00000003_sig0000040b : STD_LOGIC; 
  signal blk00000003_sig0000040a : STD_LOGIC; 
  signal blk00000003_sig00000409 : STD_LOGIC; 
  signal blk00000003_sig00000408 : STD_LOGIC; 
  signal blk00000003_sig00000407 : STD_LOGIC; 
  signal blk00000003_sig00000406 : STD_LOGIC; 
  signal blk00000003_sig00000405 : STD_LOGIC; 
  signal blk00000003_sig00000404 : STD_LOGIC; 
  signal blk00000003_sig00000403 : STD_LOGIC; 
  signal blk00000003_sig00000402 : STD_LOGIC; 
  signal blk00000003_sig00000401 : STD_LOGIC; 
  signal blk00000003_sig00000400 : STD_LOGIC; 
  signal blk00000003_sig000003ff : STD_LOGIC; 
  signal blk00000003_sig000003fe : STD_LOGIC; 
  signal blk00000003_sig000003fd : STD_LOGIC; 
  signal blk00000003_sig000003fc : STD_LOGIC; 
  signal blk00000003_sig000003fb : STD_LOGIC; 
  signal blk00000003_sig000003fa : STD_LOGIC; 
  signal blk00000003_sig000003f9 : STD_LOGIC; 
  signal blk00000003_sig000003f8 : STD_LOGIC; 
  signal blk00000003_sig000003f7 : STD_LOGIC; 
  signal blk00000003_sig000003f6 : STD_LOGIC; 
  signal blk00000003_sig000003f5 : STD_LOGIC; 
  signal blk00000003_sig000003f4 : STD_LOGIC; 
  signal blk00000003_sig000003f3 : STD_LOGIC; 
  signal blk00000003_sig000003f2 : STD_LOGIC; 
  signal blk00000003_sig000003f1 : STD_LOGIC; 
  signal blk00000003_sig000003f0 : STD_LOGIC; 
  signal blk00000003_sig000003ef : STD_LOGIC; 
  signal blk00000003_sig000003ee : STD_LOGIC; 
  signal blk00000003_sig000003ed : STD_LOGIC; 
  signal blk00000003_sig000003ec : STD_LOGIC; 
  signal blk00000003_sig000003eb : STD_LOGIC; 
  signal blk00000003_sig000003ea : STD_LOGIC; 
  signal blk00000003_sig000003e9 : STD_LOGIC; 
  signal blk00000003_sig000003e8 : STD_LOGIC; 
  signal blk00000003_sig000003e7 : STD_LOGIC; 
  signal blk00000003_sig000003e6 : STD_LOGIC; 
  signal blk00000003_sig000003e5 : STD_LOGIC; 
  signal blk00000003_sig000003e4 : STD_LOGIC; 
  signal blk00000003_sig000003e3 : STD_LOGIC; 
  signal blk00000003_sig000003e2 : STD_LOGIC; 
  signal blk00000003_sig000003e1 : STD_LOGIC; 
  signal blk00000003_sig000003e0 : STD_LOGIC; 
  signal blk00000003_sig000003df : STD_LOGIC; 
  signal blk00000003_sig000003de : STD_LOGIC; 
  signal blk00000003_sig000003dd : STD_LOGIC; 
  signal blk00000003_sig000003dc : STD_LOGIC; 
  signal blk00000003_sig000003db : STD_LOGIC; 
  signal blk00000003_sig000003da : STD_LOGIC; 
  signal blk00000003_sig000003d9 : STD_LOGIC; 
  signal blk00000003_sig000003d8 : STD_LOGIC; 
  signal blk00000003_sig000003d7 : STD_LOGIC; 
  signal blk00000003_sig000003d6 : STD_LOGIC; 
  signal blk00000003_sig000003d5 : STD_LOGIC; 
  signal blk00000003_sig000003d4 : STD_LOGIC; 
  signal blk00000003_sig000003d3 : STD_LOGIC; 
  signal blk00000003_sig000003d2 : STD_LOGIC; 
  signal blk00000003_sig000003d1 : STD_LOGIC; 
  signal blk00000003_sig000003d0 : STD_LOGIC; 
  signal blk00000003_sig000003cf : STD_LOGIC; 
  signal blk00000003_sig000003ce : STD_LOGIC; 
  signal blk00000003_sig000003cd : STD_LOGIC; 
  signal blk00000003_sig000003cc : STD_LOGIC; 
  signal blk00000003_sig000003cb : STD_LOGIC; 
  signal blk00000003_sig000003ca : STD_LOGIC; 
  signal blk00000003_sig000003c9 : STD_LOGIC; 
  signal blk00000003_sig000003c8 : STD_LOGIC; 
  signal blk00000003_sig000003c7 : STD_LOGIC; 
  signal blk00000003_sig000003c6 : STD_LOGIC; 
  signal blk00000003_sig000003c5 : STD_LOGIC; 
  signal blk00000003_sig000003c4 : STD_LOGIC; 
  signal blk00000003_sig000003c3 : STD_LOGIC; 
  signal blk00000003_sig000003c2 : STD_LOGIC; 
  signal blk00000003_sig000003c1 : STD_LOGIC; 
  signal blk00000003_sig000003c0 : STD_LOGIC; 
  signal blk00000003_sig000003bf : STD_LOGIC; 
  signal blk00000003_sig000003be : STD_LOGIC; 
  signal blk00000003_sig000003bd : STD_LOGIC; 
  signal blk00000003_sig000003bc : STD_LOGIC; 
  signal blk00000003_sig000003bb : STD_LOGIC; 
  signal blk00000003_sig000003ba : STD_LOGIC; 
  signal blk00000003_sig000003b9 : STD_LOGIC; 
  signal blk00000003_sig000003b8 : STD_LOGIC; 
  signal blk00000003_sig000003b7 : STD_LOGIC; 
  signal blk00000003_sig000003b6 : STD_LOGIC; 
  signal blk00000003_sig000003b5 : STD_LOGIC; 
  signal blk00000003_sig000003b4 : STD_LOGIC; 
  signal blk00000003_sig000003b3 : STD_LOGIC; 
  signal blk00000003_sig000003b2 : STD_LOGIC; 
  signal blk00000003_sig000003b1 : STD_LOGIC; 
  signal blk00000003_sig000003b0 : STD_LOGIC; 
  signal blk00000003_sig000003af : STD_LOGIC; 
  signal blk00000003_sig000003ae : STD_LOGIC; 
  signal blk00000003_sig000003ad : STD_LOGIC; 
  signal blk00000003_sig000003ac : STD_LOGIC; 
  signal blk00000003_sig000003ab : STD_LOGIC; 
  signal blk00000003_sig000003aa : STD_LOGIC; 
  signal blk00000003_sig000003a9 : STD_LOGIC; 
  signal blk00000003_sig000003a8 : STD_LOGIC; 
  signal blk00000003_sig000003a7 : STD_LOGIC; 
  signal blk00000003_sig000003a6 : STD_LOGIC; 
  signal blk00000003_sig000003a5 : STD_LOGIC; 
  signal blk00000003_sig000003a4 : STD_LOGIC; 
  signal blk00000003_sig000003a3 : STD_LOGIC; 
  signal blk00000003_sig000003a2 : STD_LOGIC; 
  signal blk00000003_sig000003a1 : STD_LOGIC; 
  signal blk00000003_sig000003a0 : STD_LOGIC; 
  signal blk00000003_sig0000039f : STD_LOGIC; 
  signal blk00000003_sig0000039e : STD_LOGIC; 
  signal blk00000003_sig0000039d : STD_LOGIC; 
  signal blk00000003_sig0000039c : STD_LOGIC; 
  signal blk00000003_sig0000039b : STD_LOGIC; 
  signal blk00000003_sig0000039a : STD_LOGIC; 
  signal blk00000003_sig00000399 : STD_LOGIC; 
  signal blk00000003_sig00000398 : STD_LOGIC; 
  signal blk00000003_sig00000397 : STD_LOGIC; 
  signal blk00000003_sig00000396 : STD_LOGIC; 
  signal blk00000003_sig00000395 : STD_LOGIC; 
  signal blk00000003_sig00000394 : STD_LOGIC; 
  signal blk00000003_sig00000393 : STD_LOGIC; 
  signal blk00000003_sig00000392 : STD_LOGIC; 
  signal blk00000003_sig00000391 : STD_LOGIC; 
  signal blk00000003_sig00000390 : STD_LOGIC; 
  signal blk00000003_sig0000038f : STD_LOGIC; 
  signal blk00000003_sig0000038e : STD_LOGIC; 
  signal blk00000003_sig0000038d : STD_LOGIC; 
  signal blk00000003_sig0000038c : STD_LOGIC; 
  signal blk00000003_sig0000038b : STD_LOGIC; 
  signal blk00000003_sig0000038a : STD_LOGIC; 
  signal blk00000003_sig00000389 : STD_LOGIC; 
  signal blk00000003_sig00000388 : STD_LOGIC; 
  signal blk00000003_sig00000387 : STD_LOGIC; 
  signal blk00000003_sig00000386 : STD_LOGIC; 
  signal blk00000003_sig00000385 : STD_LOGIC; 
  signal blk00000003_sig00000384 : STD_LOGIC; 
  signal blk00000003_sig00000383 : STD_LOGIC; 
  signal blk00000003_sig00000382 : STD_LOGIC; 
  signal blk00000003_sig00000381 : STD_LOGIC; 
  signal blk00000003_sig00000380 : STD_LOGIC; 
  signal blk00000003_sig0000037f : STD_LOGIC; 
  signal blk00000003_sig0000037e : STD_LOGIC; 
  signal blk00000003_sig0000037d : STD_LOGIC; 
  signal blk00000003_sig0000037c : STD_LOGIC; 
  signal blk00000003_sig0000037b : STD_LOGIC; 
  signal blk00000003_sig0000037a : STD_LOGIC; 
  signal blk00000003_sig00000379 : STD_LOGIC; 
  signal blk00000003_sig00000378 : STD_LOGIC; 
  signal blk00000003_sig00000377 : STD_LOGIC; 
  signal blk00000003_sig00000376 : STD_LOGIC; 
  signal blk00000003_sig00000375 : STD_LOGIC; 
  signal blk00000003_sig00000374 : STD_LOGIC; 
  signal blk00000003_sig00000373 : STD_LOGIC; 
  signal blk00000003_sig00000372 : STD_LOGIC; 
  signal blk00000003_sig00000371 : STD_LOGIC; 
  signal blk00000003_sig00000370 : STD_LOGIC; 
  signal blk00000003_sig0000036f : STD_LOGIC; 
  signal blk00000003_sig0000036e : STD_LOGIC; 
  signal blk00000003_sig0000036d : STD_LOGIC; 
  signal blk00000003_sig0000036c : STD_LOGIC; 
  signal blk00000003_sig0000036b : STD_LOGIC; 
  signal blk00000003_sig0000036a : STD_LOGIC; 
  signal blk00000003_sig00000369 : STD_LOGIC; 
  signal blk00000003_sig00000368 : STD_LOGIC; 
  signal blk00000003_sig00000367 : STD_LOGIC; 
  signal blk00000003_sig00000366 : STD_LOGIC; 
  signal blk00000003_sig00000365 : STD_LOGIC; 
  signal blk00000003_sig00000364 : STD_LOGIC; 
  signal blk00000003_sig00000363 : STD_LOGIC; 
  signal blk00000003_sig00000362 : STD_LOGIC; 
  signal blk00000003_sig00000361 : STD_LOGIC; 
  signal blk00000003_sig00000360 : STD_LOGIC; 
  signal blk00000003_sig0000035f : STD_LOGIC; 
  signal blk00000003_sig0000035e : STD_LOGIC; 
  signal blk00000003_sig0000035d : STD_LOGIC; 
  signal blk00000003_sig0000035c : STD_LOGIC; 
  signal blk00000003_sig0000035b : STD_LOGIC; 
  signal blk00000003_sig0000035a : STD_LOGIC; 
  signal blk00000003_sig00000359 : STD_LOGIC; 
  signal blk00000003_sig00000358 : STD_LOGIC; 
  signal blk00000003_sig00000357 : STD_LOGIC; 
  signal blk00000003_sig00000356 : STD_LOGIC; 
  signal blk00000003_sig00000355 : STD_LOGIC; 
  signal blk00000003_sig00000354 : STD_LOGIC; 
  signal blk00000003_sig00000353 : STD_LOGIC; 
  signal blk00000003_sig00000352 : STD_LOGIC; 
  signal blk00000003_sig00000351 : STD_LOGIC; 
  signal blk00000003_sig00000350 : STD_LOGIC; 
  signal blk00000003_sig0000034f : STD_LOGIC; 
  signal blk00000003_sig0000034e : STD_LOGIC; 
  signal blk00000003_sig0000034d : STD_LOGIC; 
  signal blk00000003_sig0000034c : STD_LOGIC; 
  signal blk00000003_sig0000034b : STD_LOGIC; 
  signal blk00000003_sig0000034a : STD_LOGIC; 
  signal blk00000003_sig00000349 : STD_LOGIC; 
  signal blk00000003_sig00000348 : STD_LOGIC; 
  signal blk00000003_sig00000347 : STD_LOGIC; 
  signal blk00000003_sig00000346 : STD_LOGIC; 
  signal blk00000003_sig00000345 : STD_LOGIC; 
  signal blk00000003_sig00000344 : STD_LOGIC; 
  signal blk00000003_sig00000343 : STD_LOGIC; 
  signal blk00000003_sig00000342 : STD_LOGIC; 
  signal blk00000003_sig00000341 : STD_LOGIC; 
  signal blk00000003_sig00000340 : STD_LOGIC; 
  signal blk00000003_sig0000033f : STD_LOGIC; 
  signal blk00000003_sig0000033e : STD_LOGIC; 
  signal blk00000003_sig0000033d : STD_LOGIC; 
  signal blk00000003_sig0000033c : STD_LOGIC; 
  signal blk00000003_sig0000033b : STD_LOGIC; 
  signal blk00000003_sig0000033a : STD_LOGIC; 
  signal blk00000003_sig00000339 : STD_LOGIC; 
  signal blk00000003_sig00000338 : STD_LOGIC; 
  signal blk00000003_sig00000337 : STD_LOGIC; 
  signal blk00000003_sig00000336 : STD_LOGIC; 
  signal blk00000003_sig00000335 : STD_LOGIC; 
  signal blk00000003_sig00000334 : STD_LOGIC; 
  signal blk00000003_sig00000333 : STD_LOGIC; 
  signal blk00000003_sig00000332 : STD_LOGIC; 
  signal blk00000003_sig00000331 : STD_LOGIC; 
  signal blk00000003_sig00000330 : STD_LOGIC; 
  signal blk00000003_sig0000032f : STD_LOGIC; 
  signal blk00000003_sig0000032e : STD_LOGIC; 
  signal blk00000003_sig0000032d : STD_LOGIC; 
  signal blk00000003_sig0000032c : STD_LOGIC; 
  signal blk00000003_sig0000032b : STD_LOGIC; 
  signal blk00000003_sig0000032a : STD_LOGIC; 
  signal blk00000003_sig00000329 : STD_LOGIC; 
  signal blk00000003_sig00000328 : STD_LOGIC; 
  signal blk00000003_sig00000327 : STD_LOGIC; 
  signal blk00000003_sig00000326 : STD_LOGIC; 
  signal blk00000003_sig00000325 : STD_LOGIC; 
  signal blk00000003_sig00000324 : STD_LOGIC; 
  signal blk00000003_sig00000323 : STD_LOGIC; 
  signal blk00000003_sig00000322 : STD_LOGIC; 
  signal blk00000003_sig00000321 : STD_LOGIC; 
  signal blk00000003_sig00000320 : STD_LOGIC; 
  signal blk00000003_sig0000031f : STD_LOGIC; 
  signal blk00000003_sig0000031e : STD_LOGIC; 
  signal blk00000003_sig0000031d : STD_LOGIC; 
  signal blk00000003_sig0000031c : STD_LOGIC; 
  signal blk00000003_sig0000031b : STD_LOGIC; 
  signal blk00000003_sig0000031a : STD_LOGIC; 
  signal blk00000003_sig00000319 : STD_LOGIC; 
  signal blk00000003_sig00000318 : STD_LOGIC; 
  signal blk00000003_sig00000317 : STD_LOGIC; 
  signal blk00000003_sig00000316 : STD_LOGIC; 
  signal blk00000003_sig00000315 : STD_LOGIC; 
  signal blk00000003_sig00000314 : STD_LOGIC; 
  signal blk00000003_sig00000313 : STD_LOGIC; 
  signal blk00000003_sig00000312 : STD_LOGIC; 
  signal blk00000003_sig00000311 : STD_LOGIC; 
  signal blk00000003_sig00000310 : STD_LOGIC; 
  signal blk00000003_sig0000030f : STD_LOGIC; 
  signal blk00000003_sig0000030e : STD_LOGIC; 
  signal blk00000003_sig0000030d : STD_LOGIC; 
  signal blk00000003_sig0000030c : STD_LOGIC; 
  signal blk00000003_sig0000030b : STD_LOGIC; 
  signal blk00000003_sig0000030a : STD_LOGIC; 
  signal blk00000003_sig00000309 : STD_LOGIC; 
  signal blk00000003_sig00000308 : STD_LOGIC; 
  signal blk00000003_sig00000307 : STD_LOGIC; 
  signal blk00000003_sig00000306 : STD_LOGIC; 
  signal blk00000003_sig00000305 : STD_LOGIC; 
  signal blk00000003_sig00000304 : STD_LOGIC; 
  signal blk00000003_sig00000303 : STD_LOGIC; 
  signal blk00000003_sig00000302 : STD_LOGIC; 
  signal blk00000003_sig00000301 : STD_LOGIC; 
  signal blk00000003_sig00000300 : STD_LOGIC; 
  signal blk00000003_sig000002ff : STD_LOGIC; 
  signal blk00000003_sig000002fe : STD_LOGIC; 
  signal blk00000003_sig000002fd : STD_LOGIC; 
  signal blk00000003_sig000002fc : STD_LOGIC; 
  signal blk00000003_sig000002fb : STD_LOGIC; 
  signal blk00000003_sig000002fa : STD_LOGIC; 
  signal blk00000003_sig000002f9 : STD_LOGIC; 
  signal blk00000003_sig000002f8 : STD_LOGIC; 
  signal blk00000003_sig000002f7 : STD_LOGIC; 
  signal blk00000003_sig000002f6 : STD_LOGIC; 
  signal blk00000003_sig000002f5 : STD_LOGIC; 
  signal blk00000003_sig000002f4 : STD_LOGIC; 
  signal blk00000003_sig000002f3 : STD_LOGIC; 
  signal blk00000003_sig000002f2 : STD_LOGIC; 
  signal blk00000003_sig000002f1 : STD_LOGIC; 
  signal blk00000003_sig000002f0 : STD_LOGIC; 
  signal blk00000003_sig000002ef : STD_LOGIC; 
  signal blk00000003_sig000002ee : STD_LOGIC; 
  signal blk00000003_sig000002ed : STD_LOGIC; 
  signal blk00000003_sig000002ec : STD_LOGIC; 
  signal blk00000003_sig000002eb : STD_LOGIC; 
  signal blk00000003_sig000002ea : STD_LOGIC; 
  signal blk00000003_sig000002e9 : STD_LOGIC; 
  signal blk00000003_sig000002e8 : STD_LOGIC; 
  signal blk00000003_sig000002e7 : STD_LOGIC; 
  signal blk00000003_sig000002e6 : STD_LOGIC; 
  signal blk00000003_sig000002e5 : STD_LOGIC; 
  signal blk00000003_sig000002e4 : STD_LOGIC; 
  signal blk00000003_sig000002e3 : STD_LOGIC; 
  signal blk00000003_sig000002e2 : STD_LOGIC; 
  signal blk00000003_sig000002e1 : STD_LOGIC; 
  signal blk00000003_sig000002e0 : STD_LOGIC; 
  signal blk00000003_sig000002df : STD_LOGIC; 
  signal blk00000003_sig000002de : STD_LOGIC; 
  signal blk00000003_sig000002dd : STD_LOGIC; 
  signal blk00000003_sig000002dc : STD_LOGIC; 
  signal blk00000003_sig000002db : STD_LOGIC; 
  signal blk00000003_sig000002da : STD_LOGIC; 
  signal blk00000003_sig000002d9 : STD_LOGIC; 
  signal blk00000003_sig000002d8 : STD_LOGIC; 
  signal blk00000003_sig000002d7 : STD_LOGIC; 
  signal blk00000003_sig000002d6 : STD_LOGIC; 
  signal blk00000003_sig000002d5 : STD_LOGIC; 
  signal blk00000003_sig000002d4 : STD_LOGIC; 
  signal blk00000003_sig000002d3 : STD_LOGIC; 
  signal blk00000003_sig000002d2 : STD_LOGIC; 
  signal blk00000003_sig000002d1 : STD_LOGIC; 
  signal blk00000003_sig000002d0 : STD_LOGIC; 
  signal blk00000003_sig000002cf : STD_LOGIC; 
  signal blk00000003_sig000002ce : STD_LOGIC; 
  signal blk00000003_sig000002cd : STD_LOGIC; 
  signal blk00000003_sig000002cc : STD_LOGIC; 
  signal blk00000003_sig000002cb : STD_LOGIC; 
  signal blk00000003_sig000002ca : STD_LOGIC; 
  signal blk00000003_sig000002c9 : STD_LOGIC; 
  signal blk00000003_sig000002c8 : STD_LOGIC; 
  signal blk00000003_sig000002c7 : STD_LOGIC; 
  signal blk00000003_sig000002c6 : STD_LOGIC; 
  signal blk00000003_sig000002c5 : STD_LOGIC; 
  signal blk00000003_sig000002c4 : STD_LOGIC; 
  signal blk00000003_sig000002c3 : STD_LOGIC; 
  signal blk00000003_sig000002c2 : STD_LOGIC; 
  signal blk00000003_sig000002c1 : STD_LOGIC; 
  signal blk00000003_sig000002c0 : STD_LOGIC; 
  signal blk00000003_sig000002bf : STD_LOGIC; 
  signal blk00000003_sig000002be : STD_LOGIC; 
  signal blk00000003_sig000002bd : STD_LOGIC; 
  signal blk00000003_sig000002bc : STD_LOGIC; 
  signal blk00000003_sig000002bb : STD_LOGIC; 
  signal blk00000003_sig000002ba : STD_LOGIC; 
  signal blk00000003_sig000002b9 : STD_LOGIC; 
  signal blk00000003_sig000002b8 : STD_LOGIC; 
  signal blk00000003_sig000002b7 : STD_LOGIC; 
  signal blk00000003_sig000002b6 : STD_LOGIC; 
  signal blk00000003_sig000002b5 : STD_LOGIC; 
  signal blk00000003_sig000002b4 : STD_LOGIC; 
  signal blk00000003_sig000002b3 : STD_LOGIC; 
  signal blk00000003_sig000002b2 : STD_LOGIC; 
  signal blk00000003_sig000002b1 : STD_LOGIC; 
  signal blk00000003_sig000002b0 : STD_LOGIC; 
  signal blk00000003_sig000002af : STD_LOGIC; 
  signal blk00000003_sig000002ae : STD_LOGIC; 
  signal blk00000003_sig000002ad : STD_LOGIC; 
  signal blk00000003_sig000002ac : STD_LOGIC; 
  signal blk00000003_sig000002ab : STD_LOGIC; 
  signal blk00000003_sig000002aa : STD_LOGIC; 
  signal blk00000003_sig000002a9 : STD_LOGIC; 
  signal blk00000003_sig000002a8 : STD_LOGIC; 
  signal blk00000003_sig000002a7 : STD_LOGIC; 
  signal blk00000003_sig000002a6 : STD_LOGIC; 
  signal blk00000003_sig000002a5 : STD_LOGIC; 
  signal blk00000003_sig000002a4 : STD_LOGIC; 
  signal blk00000003_sig000002a3 : STD_LOGIC; 
  signal blk00000003_sig000002a2 : STD_LOGIC; 
  signal blk00000003_sig000002a1 : STD_LOGIC; 
  signal blk00000003_sig000002a0 : STD_LOGIC; 
  signal blk00000003_sig0000029f : STD_LOGIC; 
  signal blk00000003_sig0000029e : STD_LOGIC; 
  signal blk00000003_sig0000029d : STD_LOGIC; 
  signal blk00000003_sig0000029c : STD_LOGIC; 
  signal blk00000003_sig0000029b : STD_LOGIC; 
  signal blk00000003_sig0000029a : STD_LOGIC; 
  signal blk00000003_sig00000299 : STD_LOGIC; 
  signal blk00000003_sig00000298 : STD_LOGIC; 
  signal blk00000003_sig00000297 : STD_LOGIC; 
  signal blk00000003_sig00000296 : STD_LOGIC; 
  signal blk00000003_sig00000295 : STD_LOGIC; 
  signal blk00000003_sig00000294 : STD_LOGIC; 
  signal blk00000003_sig00000293 : STD_LOGIC; 
  signal blk00000003_sig00000292 : STD_LOGIC; 
  signal blk00000003_sig00000291 : STD_LOGIC; 
  signal blk00000003_sig00000290 : STD_LOGIC; 
  signal blk00000003_sig0000028f : STD_LOGIC; 
  signal blk00000003_sig0000028e : STD_LOGIC; 
  signal blk00000003_sig0000028d : STD_LOGIC; 
  signal blk00000003_sig0000028c : STD_LOGIC; 
  signal blk00000003_sig0000028b : STD_LOGIC; 
  signal blk00000003_sig0000028a : STD_LOGIC; 
  signal blk00000003_sig00000289 : STD_LOGIC; 
  signal blk00000003_sig00000288 : STD_LOGIC; 
  signal blk00000003_sig00000287 : STD_LOGIC; 
  signal blk00000003_sig00000286 : STD_LOGIC; 
  signal blk00000003_sig00000285 : STD_LOGIC; 
  signal blk00000003_sig00000284 : STD_LOGIC; 
  signal blk00000003_sig00000283 : STD_LOGIC; 
  signal blk00000003_sig00000282 : STD_LOGIC; 
  signal blk00000003_sig00000281 : STD_LOGIC; 
  signal blk00000003_sig00000280 : STD_LOGIC; 
  signal blk00000003_sig0000027f : STD_LOGIC; 
  signal blk00000003_sig0000027e : STD_LOGIC; 
  signal blk00000003_sig0000027d : STD_LOGIC; 
  signal blk00000003_sig0000027c : STD_LOGIC; 
  signal blk00000003_sig0000027b : STD_LOGIC; 
  signal blk00000003_sig0000027a : STD_LOGIC; 
  signal blk00000003_sig00000279 : STD_LOGIC; 
  signal blk00000003_sig00000278 : STD_LOGIC; 
  signal blk00000003_sig00000277 : STD_LOGIC; 
  signal blk00000003_sig00000276 : STD_LOGIC; 
  signal blk00000003_sig00000275 : STD_LOGIC; 
  signal blk00000003_sig00000274 : STD_LOGIC; 
  signal blk00000003_sig00000273 : STD_LOGIC; 
  signal blk00000003_sig00000272 : STD_LOGIC; 
  signal blk00000003_sig00000271 : STD_LOGIC; 
  signal blk00000003_sig00000270 : STD_LOGIC; 
  signal blk00000003_sig0000026f : STD_LOGIC; 
  signal blk00000003_sig0000026e : STD_LOGIC; 
  signal blk00000003_sig0000026d : STD_LOGIC; 
  signal blk00000003_sig0000026c : STD_LOGIC; 
  signal blk00000003_sig0000026b : STD_LOGIC; 
  signal blk00000003_sig0000026a : STD_LOGIC; 
  signal blk00000003_sig00000269 : STD_LOGIC; 
  signal blk00000003_sig00000268 : STD_LOGIC; 
  signal blk00000003_sig00000267 : STD_LOGIC; 
  signal blk00000003_sig00000266 : STD_LOGIC; 
  signal blk00000003_sig00000265 : STD_LOGIC; 
  signal blk00000003_sig00000264 : STD_LOGIC; 
  signal blk00000003_sig00000263 : STD_LOGIC; 
  signal blk00000003_sig00000262 : STD_LOGIC; 
  signal blk00000003_sig00000261 : STD_LOGIC; 
  signal blk00000003_sig00000260 : STD_LOGIC; 
  signal blk00000003_sig0000025f : STD_LOGIC; 
  signal blk00000003_sig0000025e : STD_LOGIC; 
  signal blk00000003_sig0000025d : STD_LOGIC; 
  signal blk00000003_sig0000025c : STD_LOGIC; 
  signal blk00000003_sig0000025b : STD_LOGIC; 
  signal blk00000003_sig0000025a : STD_LOGIC; 
  signal blk00000003_sig00000259 : STD_LOGIC; 
  signal blk00000003_sig00000258 : STD_LOGIC; 
  signal blk00000003_sig00000257 : STD_LOGIC; 
  signal blk00000003_sig00000256 : STD_LOGIC; 
  signal blk00000003_sig00000255 : STD_LOGIC; 
  signal blk00000003_sig00000254 : STD_LOGIC; 
  signal blk00000003_sig00000253 : STD_LOGIC; 
  signal blk00000003_sig00000252 : STD_LOGIC; 
  signal blk00000003_sig00000251 : STD_LOGIC; 
  signal blk00000003_sig00000250 : STD_LOGIC; 
  signal blk00000003_sig0000024f : STD_LOGIC; 
  signal blk00000003_sig0000024e : STD_LOGIC; 
  signal blk00000003_sig0000024d : STD_LOGIC; 
  signal blk00000003_sig0000024c : STD_LOGIC; 
  signal blk00000003_sig0000024b : STD_LOGIC; 
  signal blk00000003_sig0000024a : STD_LOGIC; 
  signal blk00000003_sig00000249 : STD_LOGIC; 
  signal blk00000003_sig00000248 : STD_LOGIC; 
  signal blk00000003_sig00000247 : STD_LOGIC; 
  signal blk00000003_sig00000246 : STD_LOGIC; 
  signal blk00000003_sig00000245 : STD_LOGIC; 
  signal blk00000003_sig00000244 : STD_LOGIC; 
  signal blk00000003_sig00000243 : STD_LOGIC; 
  signal blk00000003_sig00000242 : STD_LOGIC; 
  signal blk00000003_sig00000241 : STD_LOGIC; 
  signal blk00000003_sig00000240 : STD_LOGIC; 
  signal blk00000003_sig0000023f : STD_LOGIC; 
  signal blk00000003_sig0000023e : STD_LOGIC; 
  signal blk00000003_sig0000023d : STD_LOGIC; 
  signal blk00000003_sig0000023c : STD_LOGIC; 
  signal blk00000003_sig0000023b : STD_LOGIC; 
  signal blk00000003_sig0000023a : STD_LOGIC; 
  signal blk00000003_sig00000239 : STD_LOGIC; 
  signal blk00000003_sig00000238 : STD_LOGIC; 
  signal blk00000003_sig00000237 : STD_LOGIC; 
  signal blk00000003_sig00000236 : STD_LOGIC; 
  signal blk00000003_sig00000235 : STD_LOGIC; 
  signal blk00000003_sig00000234 : STD_LOGIC; 
  signal blk00000003_sig00000233 : STD_LOGIC; 
  signal blk00000003_sig00000232 : STD_LOGIC; 
  signal blk00000003_sig00000231 : STD_LOGIC; 
  signal blk00000003_sig00000230 : STD_LOGIC; 
  signal blk00000003_sig0000022f : STD_LOGIC; 
  signal blk00000003_sig0000022e : STD_LOGIC; 
  signal blk00000003_sig0000022d : STD_LOGIC; 
  signal blk00000003_sig0000022c : STD_LOGIC; 
  signal blk00000003_sig0000022b : STD_LOGIC; 
  signal blk00000003_sig0000022a : STD_LOGIC; 
  signal blk00000003_sig00000229 : STD_LOGIC; 
  signal blk00000003_sig00000228 : STD_LOGIC; 
  signal blk00000003_sig00000227 : STD_LOGIC; 
  signal blk00000003_sig00000226 : STD_LOGIC; 
  signal blk00000003_sig00000225 : STD_LOGIC; 
  signal blk00000003_sig00000224 : STD_LOGIC; 
  signal blk00000003_sig00000223 : STD_LOGIC; 
  signal blk00000003_sig00000222 : STD_LOGIC; 
  signal blk00000003_sig00000221 : STD_LOGIC; 
  signal blk00000003_sig00000220 : STD_LOGIC; 
  signal blk00000003_sig0000021f : STD_LOGIC; 
  signal blk00000003_sig0000021e : STD_LOGIC; 
  signal blk00000003_sig0000021d : STD_LOGIC; 
  signal blk00000003_sig0000021c : STD_LOGIC; 
  signal blk00000003_sig0000021b : STD_LOGIC; 
  signal blk00000003_sig0000021a : STD_LOGIC; 
  signal blk00000003_sig00000219 : STD_LOGIC; 
  signal blk00000003_sig00000218 : STD_LOGIC; 
  signal blk00000003_sig00000217 : STD_LOGIC; 
  signal blk00000003_sig00000216 : STD_LOGIC; 
  signal blk00000003_sig00000215 : STD_LOGIC; 
  signal blk00000003_sig00000214 : STD_LOGIC; 
  signal blk00000003_sig00000213 : STD_LOGIC; 
  signal blk00000003_sig00000212 : STD_LOGIC; 
  signal blk00000003_sig00000211 : STD_LOGIC; 
  signal blk00000003_sig00000210 : STD_LOGIC; 
  signal blk00000003_sig0000020f : STD_LOGIC; 
  signal blk00000003_sig0000020e : STD_LOGIC; 
  signal blk00000003_sig0000020d : STD_LOGIC; 
  signal blk00000003_sig0000020c : STD_LOGIC; 
  signal blk00000003_sig0000020b : STD_LOGIC; 
  signal blk00000003_sig0000020a : STD_LOGIC; 
  signal blk00000003_sig00000209 : STD_LOGIC; 
  signal blk00000003_sig00000208 : STD_LOGIC; 
  signal blk00000003_sig00000207 : STD_LOGIC; 
  signal blk00000003_sig00000206 : STD_LOGIC; 
  signal blk00000003_sig00000205 : STD_LOGIC; 
  signal blk00000003_sig00000204 : STD_LOGIC; 
  signal blk00000003_sig00000203 : STD_LOGIC; 
  signal blk00000003_sig00000202 : STD_LOGIC; 
  signal blk00000003_sig00000201 : STD_LOGIC; 
  signal blk00000003_sig00000200 : STD_LOGIC; 
  signal blk00000003_sig000001ff : STD_LOGIC; 
  signal blk00000003_sig000001fe : STD_LOGIC; 
  signal blk00000003_sig000001fd : STD_LOGIC; 
  signal blk00000003_sig000001fc : STD_LOGIC; 
  signal blk00000003_sig000001fb : STD_LOGIC; 
  signal blk00000003_sig000001fa : STD_LOGIC; 
  signal blk00000003_sig000001f9 : STD_LOGIC; 
  signal blk00000003_sig000001f8 : STD_LOGIC; 
  signal blk00000003_sig000001f7 : STD_LOGIC; 
  signal blk00000003_sig000001f6 : STD_LOGIC; 
  signal blk00000003_sig000001f5 : STD_LOGIC; 
  signal blk00000003_sig000001f4 : STD_LOGIC; 
  signal blk00000003_sig000001f3 : STD_LOGIC; 
  signal blk00000003_sig000001f2 : STD_LOGIC; 
  signal blk00000003_sig000001f1 : STD_LOGIC; 
  signal blk00000003_sig000001f0 : STD_LOGIC; 
  signal blk00000003_sig000001ef : STD_LOGIC; 
  signal blk00000003_sig000001ee : STD_LOGIC; 
  signal blk00000003_sig000001ed : STD_LOGIC; 
  signal blk00000003_sig000001ec : STD_LOGIC; 
  signal blk00000003_sig000001eb : STD_LOGIC; 
  signal blk00000003_sig000001ea : STD_LOGIC; 
  signal blk00000003_sig000001e9 : STD_LOGIC; 
  signal blk00000003_sig000001e8 : STD_LOGIC; 
  signal blk00000003_sig000001e7 : STD_LOGIC; 
  signal blk00000003_sig000001e6 : STD_LOGIC; 
  signal blk00000003_sig000001e5 : STD_LOGIC; 
  signal blk00000003_sig000001e4 : STD_LOGIC; 
  signal blk00000003_sig000001e3 : STD_LOGIC; 
  signal blk00000003_sig000001e2 : STD_LOGIC; 
  signal blk00000003_sig000001e1 : STD_LOGIC; 
  signal blk00000003_sig000001e0 : STD_LOGIC; 
  signal blk00000003_sig000001df : STD_LOGIC; 
  signal blk00000003_sig000001de : STD_LOGIC; 
  signal blk00000003_sig000001dd : STD_LOGIC; 
  signal blk00000003_sig000001dc : STD_LOGIC; 
  signal blk00000003_sig000001db : STD_LOGIC; 
  signal blk00000003_sig000001da : STD_LOGIC; 
  signal blk00000003_sig000001d9 : STD_LOGIC; 
  signal blk00000003_sig000001d8 : STD_LOGIC; 
  signal blk00000003_sig000001d7 : STD_LOGIC; 
  signal blk00000003_sig000001d6 : STD_LOGIC; 
  signal blk00000003_sig000001d5 : STD_LOGIC; 
  signal blk00000003_sig000001d4 : STD_LOGIC; 
  signal blk00000003_sig000001d3 : STD_LOGIC; 
  signal blk00000003_sig000001d2 : STD_LOGIC; 
  signal blk00000003_sig000001d1 : STD_LOGIC; 
  signal blk00000003_sig000001d0 : STD_LOGIC; 
  signal blk00000003_sig000001cf : STD_LOGIC; 
  signal blk00000003_sig000001ce : STD_LOGIC; 
  signal blk00000003_sig000001cd : STD_LOGIC; 
  signal blk00000003_sig000001cc : STD_LOGIC; 
  signal blk00000003_sig000001cb : STD_LOGIC; 
  signal blk00000003_sig000001ca : STD_LOGIC; 
  signal blk00000003_sig000001c9 : STD_LOGIC; 
  signal blk00000003_sig000001c8 : STD_LOGIC; 
  signal blk00000003_sig000001c7 : STD_LOGIC; 
  signal blk00000003_sig000001c6 : STD_LOGIC; 
  signal blk00000003_sig000001c5 : STD_LOGIC; 
  signal blk00000003_sig000001c4 : STD_LOGIC; 
  signal blk00000003_sig000001c3 : STD_LOGIC; 
  signal blk00000003_sig000001c2 : STD_LOGIC; 
  signal blk00000003_sig000001c1 : STD_LOGIC; 
  signal blk00000003_sig000001c0 : STD_LOGIC; 
  signal blk00000003_sig000001bf : STD_LOGIC; 
  signal blk00000003_sig000001be : STD_LOGIC; 
  signal blk00000003_sig000001bd : STD_LOGIC; 
  signal blk00000003_sig000001bc : STD_LOGIC; 
  signal blk00000003_sig000001bb : STD_LOGIC; 
  signal blk00000003_sig000001ba : STD_LOGIC; 
  signal blk00000003_sig000001b9 : STD_LOGIC; 
  signal blk00000003_sig000001b8 : STD_LOGIC; 
  signal blk00000003_sig000001b7 : STD_LOGIC; 
  signal blk00000003_sig000001b6 : STD_LOGIC; 
  signal blk00000003_sig000001b5 : STD_LOGIC; 
  signal blk00000003_sig000001b4 : STD_LOGIC; 
  signal blk00000003_sig000001b3 : STD_LOGIC; 
  signal blk00000003_sig000001b2 : STD_LOGIC; 
  signal blk00000003_sig000001b1 : STD_LOGIC; 
  signal blk00000003_sig000001b0 : STD_LOGIC; 
  signal blk00000003_sig000001af : STD_LOGIC; 
  signal blk00000003_sig000001ae : STD_LOGIC; 
  signal blk00000003_sig000001ad : STD_LOGIC; 
  signal blk00000003_sig000001ac : STD_LOGIC; 
  signal blk00000003_sig000001ab : STD_LOGIC; 
  signal blk00000003_sig000001aa : STD_LOGIC; 
  signal blk00000003_sig000001a9 : STD_LOGIC; 
  signal blk00000003_sig000001a8 : STD_LOGIC; 
  signal blk00000003_sig000001a7 : STD_LOGIC; 
  signal blk00000003_sig000001a6 : STD_LOGIC; 
  signal blk00000003_sig000001a5 : STD_LOGIC; 
  signal blk00000003_sig000001a4 : STD_LOGIC; 
  signal blk00000003_sig000001a3 : STD_LOGIC; 
  signal blk00000003_sig000001a2 : STD_LOGIC; 
  signal blk00000003_sig000001a1 : STD_LOGIC; 
  signal blk00000003_sig000001a0 : STD_LOGIC; 
  signal blk00000003_sig0000019f : STD_LOGIC; 
  signal blk00000003_sig0000019e : STD_LOGIC; 
  signal blk00000003_sig0000019d : STD_LOGIC; 
  signal blk00000003_sig0000019c : STD_LOGIC; 
  signal blk00000003_sig0000019b : STD_LOGIC; 
  signal blk00000003_sig0000019a : STD_LOGIC; 
  signal blk00000003_sig00000199 : STD_LOGIC; 
  signal blk00000003_sig00000198 : STD_LOGIC; 
  signal blk00000003_sig00000197 : STD_LOGIC; 
  signal blk00000003_sig00000196 : STD_LOGIC; 
  signal blk00000003_sig00000195 : STD_LOGIC; 
  signal blk00000003_sig00000194 : STD_LOGIC; 
  signal blk00000003_sig00000193 : STD_LOGIC; 
  signal blk00000003_sig00000192 : STD_LOGIC; 
  signal blk00000003_sig00000191 : STD_LOGIC; 
  signal blk00000003_sig00000190 : STD_LOGIC; 
  signal blk00000003_sig0000018f : STD_LOGIC; 
  signal blk00000003_sig0000018e : STD_LOGIC; 
  signal blk00000003_sig0000018d : STD_LOGIC; 
  signal blk00000003_sig0000018c : STD_LOGIC; 
  signal blk00000003_sig0000018b : STD_LOGIC; 
  signal blk00000003_sig0000018a : STD_LOGIC; 
  signal blk00000003_sig00000189 : STD_LOGIC; 
  signal blk00000003_sig00000188 : STD_LOGIC; 
  signal blk00000003_sig00000187 : STD_LOGIC; 
  signal blk00000003_sig00000186 : STD_LOGIC; 
  signal blk00000003_sig00000185 : STD_LOGIC; 
  signal blk00000003_sig00000184 : STD_LOGIC; 
  signal blk00000003_sig00000183 : STD_LOGIC; 
  signal blk00000003_sig00000182 : STD_LOGIC; 
  signal blk00000003_sig00000181 : STD_LOGIC; 
  signal blk00000003_sig00000180 : STD_LOGIC; 
  signal blk00000003_sig0000017f : STD_LOGIC; 
  signal blk00000003_sig0000017e : STD_LOGIC; 
  signal blk00000003_sig0000017d : STD_LOGIC; 
  signal blk00000003_sig0000017c : STD_LOGIC; 
  signal blk00000003_sig0000017b : STD_LOGIC; 
  signal blk00000003_sig0000017a : STD_LOGIC; 
  signal blk00000003_sig00000179 : STD_LOGIC; 
  signal blk00000003_sig00000178 : STD_LOGIC; 
  signal blk00000003_sig00000177 : STD_LOGIC; 
  signal blk00000003_sig00000176 : STD_LOGIC; 
  signal blk00000003_sig00000175 : STD_LOGIC; 
  signal blk00000003_sig00000174 : STD_LOGIC; 
  signal blk00000003_sig00000173 : STD_LOGIC; 
  signal blk00000003_sig00000172 : STD_LOGIC; 
  signal blk00000003_sig00000171 : STD_LOGIC; 
  signal blk00000003_sig00000170 : STD_LOGIC; 
  signal blk00000003_sig0000016f : STD_LOGIC; 
  signal blk00000003_sig0000016e : STD_LOGIC; 
  signal blk00000003_sig0000016d : STD_LOGIC; 
  signal blk00000003_sig0000016c : STD_LOGIC; 
  signal blk00000003_sig0000016b : STD_LOGIC; 
  signal blk00000003_sig0000016a : STD_LOGIC; 
  signal blk00000003_sig00000169 : STD_LOGIC; 
  signal blk00000003_sig00000168 : STD_LOGIC; 
  signal blk00000003_sig00000167 : STD_LOGIC; 
  signal blk00000003_sig00000166 : STD_LOGIC; 
  signal blk00000003_sig00000165 : STD_LOGIC; 
  signal blk00000003_sig00000164 : STD_LOGIC; 
  signal blk00000003_sig00000163 : STD_LOGIC; 
  signal blk00000003_sig00000162 : STD_LOGIC; 
  signal blk00000003_sig00000161 : STD_LOGIC; 
  signal blk00000003_sig00000160 : STD_LOGIC; 
  signal blk00000003_sig0000015f : STD_LOGIC; 
  signal blk00000003_sig0000015e : STD_LOGIC; 
  signal blk00000003_sig0000015d : STD_LOGIC; 
  signal blk00000003_sig0000015c : STD_LOGIC; 
  signal blk00000003_sig0000015b : STD_LOGIC; 
  signal blk00000003_sig0000015a : STD_LOGIC; 
  signal blk00000003_sig00000159 : STD_LOGIC; 
  signal blk00000003_sig00000158 : STD_LOGIC; 
  signal blk00000003_sig00000157 : STD_LOGIC; 
  signal blk00000003_sig00000156 : STD_LOGIC; 
  signal blk00000003_sig00000155 : STD_LOGIC; 
  signal blk00000003_sig00000154 : STD_LOGIC; 
  signal blk00000003_sig00000153 : STD_LOGIC; 
  signal blk00000003_sig00000152 : STD_LOGIC; 
  signal blk00000003_sig00000151 : STD_LOGIC; 
  signal blk00000003_sig00000150 : STD_LOGIC; 
  signal blk00000003_sig0000014f : STD_LOGIC; 
  signal blk00000003_sig0000014e : STD_LOGIC; 
  signal blk00000003_sig0000014d : STD_LOGIC; 
  signal blk00000003_sig0000014c : STD_LOGIC; 
  signal blk00000003_sig0000014b : STD_LOGIC; 
  signal blk00000003_sig0000014a : STD_LOGIC; 
  signal blk00000003_sig00000149 : STD_LOGIC; 
  signal blk00000003_sig00000148 : STD_LOGIC; 
  signal blk00000003_sig00000147 : STD_LOGIC; 
  signal blk00000003_sig00000146 : STD_LOGIC; 
  signal blk00000003_sig00000145 : STD_LOGIC; 
  signal blk00000003_sig00000144 : STD_LOGIC; 
  signal blk00000003_sig00000143 : STD_LOGIC; 
  signal blk00000003_sig00000142 : STD_LOGIC; 
  signal blk00000003_sig00000141 : STD_LOGIC; 
  signal blk00000003_sig00000140 : STD_LOGIC; 
  signal blk00000003_sig0000013f : STD_LOGIC; 
  signal blk00000003_sig0000013e : STD_LOGIC; 
  signal blk00000003_sig0000013d : STD_LOGIC; 
  signal blk00000003_sig0000013c : STD_LOGIC; 
  signal blk00000003_sig0000013b : STD_LOGIC; 
  signal blk00000003_sig0000013a : STD_LOGIC; 
  signal blk00000003_sig00000139 : STD_LOGIC; 
  signal blk00000003_sig00000138 : STD_LOGIC; 
  signal blk00000003_sig00000137 : STD_LOGIC; 
  signal blk00000003_sig00000136 : STD_LOGIC; 
  signal blk00000003_sig00000135 : STD_LOGIC; 
  signal blk00000003_sig00000134 : STD_LOGIC; 
  signal blk00000003_sig00000133 : STD_LOGIC; 
  signal blk00000003_sig00000132 : STD_LOGIC; 
  signal blk00000003_sig00000131 : STD_LOGIC; 
  signal blk00000003_sig00000130 : STD_LOGIC; 
  signal blk00000003_sig0000012f : STD_LOGIC; 
  signal blk00000003_sig0000012e : STD_LOGIC; 
  signal blk00000003_sig0000012d : STD_LOGIC; 
  signal blk00000003_sig0000012c : STD_LOGIC; 
  signal blk00000003_sig0000012b : STD_LOGIC; 
  signal blk00000003_sig0000012a : STD_LOGIC; 
  signal blk00000003_sig00000129 : STD_LOGIC; 
  signal blk00000003_sig00000128 : STD_LOGIC; 
  signal blk00000003_sig00000127 : STD_LOGIC; 
  signal blk00000003_sig00000126 : STD_LOGIC; 
  signal blk00000003_sig00000125 : STD_LOGIC; 
  signal blk00000003_sig00000124 : STD_LOGIC; 
  signal blk00000003_sig00000123 : STD_LOGIC; 
  signal blk00000003_sig00000122 : STD_LOGIC; 
  signal blk00000003_sig00000121 : STD_LOGIC; 
  signal blk00000003_sig00000120 : STD_LOGIC; 
  signal blk00000003_sig0000011f : STD_LOGIC; 
  signal blk00000003_sig0000011e : STD_LOGIC; 
  signal blk00000003_sig0000011d : STD_LOGIC; 
  signal blk00000003_sig0000011c : STD_LOGIC; 
  signal blk00000003_sig0000011b : STD_LOGIC; 
  signal blk00000003_sig0000011a : STD_LOGIC; 
  signal blk00000003_sig00000119 : STD_LOGIC; 
  signal blk00000003_sig00000118 : STD_LOGIC; 
  signal blk00000003_sig00000117 : STD_LOGIC; 
  signal blk00000003_sig00000116 : STD_LOGIC; 
  signal blk00000003_sig00000115 : STD_LOGIC; 
  signal blk00000003_sig00000114 : STD_LOGIC; 
  signal blk00000003_sig00000113 : STD_LOGIC; 
  signal blk00000003_sig00000112 : STD_LOGIC; 
  signal blk00000003_sig00000111 : STD_LOGIC; 
  signal blk00000003_sig00000110 : STD_LOGIC; 
  signal blk00000003_sig0000010f : STD_LOGIC; 
  signal blk00000003_sig0000010e : STD_LOGIC; 
  signal blk00000003_sig0000010d : STD_LOGIC; 
  signal blk00000003_sig0000010c : STD_LOGIC; 
  signal blk00000003_sig0000010b : STD_LOGIC; 
  signal blk00000003_sig0000010a : STD_LOGIC; 
  signal blk00000003_sig00000109 : STD_LOGIC; 
  signal blk00000003_sig00000108 : STD_LOGIC; 
  signal blk00000003_sig00000107 : STD_LOGIC; 
  signal blk00000003_sig00000106 : STD_LOGIC; 
  signal blk00000003_sig00000105 : STD_LOGIC; 
  signal blk00000003_sig00000104 : STD_LOGIC; 
  signal blk00000003_sig00000103 : STD_LOGIC; 
  signal blk00000003_sig00000102 : STD_LOGIC; 
  signal blk00000003_sig00000101 : STD_LOGIC; 
  signal blk00000003_sig00000100 : STD_LOGIC; 
  signal blk00000003_sig000000ff : STD_LOGIC; 
  signal blk00000003_sig000000fe : STD_LOGIC; 
  signal blk00000003_sig000000fd : STD_LOGIC; 
  signal blk00000003_sig000000fc : STD_LOGIC; 
  signal blk00000003_sig000000fb : STD_LOGIC; 
  signal blk00000003_sig000000fa : STD_LOGIC; 
  signal blk00000003_sig000000f9 : STD_LOGIC; 
  signal blk00000003_sig000000f8 : STD_LOGIC; 
  signal blk00000003_sig000000f7 : STD_LOGIC; 
  signal blk00000003_sig000000f6 : STD_LOGIC; 
  signal blk00000003_sig000000f5 : STD_LOGIC; 
  signal blk00000003_sig000000f4 : STD_LOGIC; 
  signal blk00000003_sig000000f3 : STD_LOGIC; 
  signal blk00000003_sig000000f2 : STD_LOGIC; 
  signal blk00000003_sig000000f1 : STD_LOGIC; 
  signal blk00000003_sig000000f0 : STD_LOGIC; 
  signal blk00000003_sig000000ef : STD_LOGIC; 
  signal blk00000003_sig000000ee : STD_LOGIC; 
  signal blk00000003_sig000000ed : STD_LOGIC; 
  signal blk00000003_sig000000ec : STD_LOGIC; 
  signal blk00000003_sig000000eb : STD_LOGIC; 
  signal blk00000003_sig000000ea : STD_LOGIC; 
  signal blk00000003_sig000000e9 : STD_LOGIC; 
  signal blk00000003_sig000000e8 : STD_LOGIC; 
  signal blk00000003_sig000000e7 : STD_LOGIC; 
  signal blk00000003_sig000000e6 : STD_LOGIC; 
  signal blk00000003_sig000000e5 : STD_LOGIC; 
  signal blk00000003_sig000000e4 : STD_LOGIC; 
  signal blk00000003_sig000000e3 : STD_LOGIC; 
  signal blk00000003_sig000000e2 : STD_LOGIC; 
  signal blk00000003_sig000000e1 : STD_LOGIC; 
  signal blk00000003_sig000000e0 : STD_LOGIC; 
  signal blk00000003_sig000000df : STD_LOGIC; 
  signal blk00000003_sig000000de : STD_LOGIC; 
  signal blk00000003_sig000000dd : STD_LOGIC; 
  signal blk00000003_sig000000dc : STD_LOGIC; 
  signal blk00000003_sig000000db : STD_LOGIC; 
  signal blk00000003_sig000000da : STD_LOGIC; 
  signal blk00000003_sig000000d9 : STD_LOGIC; 
  signal blk00000003_sig000000d8 : STD_LOGIC; 
  signal blk00000003_sig000000d7 : STD_LOGIC; 
  signal blk00000003_sig000000d6 : STD_LOGIC; 
  signal blk00000003_sig000000d5 : STD_LOGIC; 
  signal blk00000003_sig000000d4 : STD_LOGIC; 
  signal blk00000003_sig000000d3 : STD_LOGIC; 
  signal blk00000003_sig000000d2 : STD_LOGIC; 
  signal blk00000003_sig000000d1 : STD_LOGIC; 
  signal blk00000003_sig000000d0 : STD_LOGIC; 
  signal blk00000003_sig000000cf : STD_LOGIC; 
  signal blk00000003_sig000000ce : STD_LOGIC; 
  signal blk00000003_sig000000cd : STD_LOGIC; 
  signal blk00000003_sig000000cc : STD_LOGIC; 
  signal blk00000003_sig000000cb : STD_LOGIC; 
  signal blk00000003_sig000000ca : STD_LOGIC; 
  signal blk00000003_sig000000c9 : STD_LOGIC; 
  signal blk00000003_sig000000c8 : STD_LOGIC; 
  signal blk00000003_sig000000c7 : STD_LOGIC; 
  signal blk00000003_sig000000c6 : STD_LOGIC; 
  signal blk00000003_sig000000c5 : STD_LOGIC; 
  signal blk00000003_sig000000c4 : STD_LOGIC; 
  signal blk00000003_sig000000c3 : STD_LOGIC; 
  signal blk00000003_sig000000c2 : STD_LOGIC; 
  signal blk00000003_sig000000c1 : STD_LOGIC; 
  signal blk00000003_sig000000c0 : STD_LOGIC; 
  signal blk00000003_sig000000bf : STD_LOGIC; 
  signal blk00000003_sig000000be : STD_LOGIC; 
  signal blk00000003_sig000000bd : STD_LOGIC; 
  signal blk00000003_sig000000bc : STD_LOGIC; 
  signal blk00000003_sig000000bb : STD_LOGIC; 
  signal blk00000003_sig000000ba : STD_LOGIC; 
  signal blk00000003_sig000000b9 : STD_LOGIC; 
  signal blk00000003_sig000000b8 : STD_LOGIC; 
  signal blk00000003_sig000000b7 : STD_LOGIC; 
  signal blk00000003_sig000000b6 : STD_LOGIC; 
  signal blk00000003_sig000000b5 : STD_LOGIC; 
  signal blk00000003_sig000000b4 : STD_LOGIC; 
  signal blk00000003_sig000000b3 : STD_LOGIC; 
  signal blk00000003_sig000000b2 : STD_LOGIC; 
  signal blk00000003_sig000000b1 : STD_LOGIC; 
  signal blk00000003_sig000000b0 : STD_LOGIC; 
  signal blk00000003_sig000000af : STD_LOGIC; 
  signal blk00000003_sig000000ae : STD_LOGIC; 
  signal blk00000003_sig000000ad : STD_LOGIC; 
  signal blk00000003_sig000000ac : STD_LOGIC; 
  signal blk00000003_sig000000ab : STD_LOGIC; 
  signal blk00000003_sig000000aa : STD_LOGIC; 
  signal blk00000003_sig000000a9 : STD_LOGIC; 
  signal blk00000003_sig000000a8 : STD_LOGIC; 
  signal blk00000003_sig000000a7 : STD_LOGIC; 
  signal blk00000003_sig000000a6 : STD_LOGIC; 
  signal blk00000003_sig000000a5 : STD_LOGIC; 
  signal blk00000003_sig000000a4 : STD_LOGIC; 
  signal blk00000003_sig000000a3 : STD_LOGIC; 
  signal blk00000003_sig000000a2 : STD_LOGIC; 
  signal blk00000003_sig000000a1 : STD_LOGIC; 
  signal blk00000003_sig000000a0 : STD_LOGIC; 
  signal blk00000003_sig0000009f : STD_LOGIC; 
  signal blk00000003_sig0000009e : STD_LOGIC; 
  signal blk00000003_sig0000009d : STD_LOGIC; 
  signal blk00000003_sig0000009c : STD_LOGIC; 
  signal blk00000003_sig0000009b : STD_LOGIC; 
  signal blk00000003_sig0000009a : STD_LOGIC; 
  signal blk00000003_sig00000099 : STD_LOGIC; 
  signal blk00000003_sig00000098 : STD_LOGIC; 
  signal blk00000003_sig00000097 : STD_LOGIC; 
  signal blk00000003_sig00000096 : STD_LOGIC; 
  signal blk00000003_sig00000095 : STD_LOGIC; 
  signal blk00000003_sig00000094 : STD_LOGIC; 
  signal blk00000003_sig00000093 : STD_LOGIC; 
  signal blk00000003_sig00000092 : STD_LOGIC; 
  signal blk00000003_sig00000091 : STD_LOGIC; 
  signal blk00000003_sig00000090 : STD_LOGIC; 
  signal blk00000003_sig0000008f : STD_LOGIC; 
  signal blk00000003_sig0000008e : STD_LOGIC; 
  signal blk00000003_sig0000008d : STD_LOGIC; 
  signal blk00000003_sig0000008c : STD_LOGIC; 
  signal blk00000003_sig0000008b : STD_LOGIC; 
  signal blk00000003_sig0000008a : STD_LOGIC; 
  signal blk00000003_sig00000089 : STD_LOGIC; 
  signal blk00000003_sig00000088 : STD_LOGIC; 
  signal blk00000003_sig00000087 : STD_LOGIC; 
  signal blk00000003_sig00000086 : STD_LOGIC; 
  signal blk00000003_sig00000085 : STD_LOGIC; 
  signal blk00000003_sig00000084 : STD_LOGIC; 
  signal blk00000003_sig00000083 : STD_LOGIC; 
  signal blk00000003_sig00000082 : STD_LOGIC; 
  signal blk00000003_sig00000081 : STD_LOGIC; 
  signal blk00000003_sig00000080 : STD_LOGIC; 
  signal blk00000003_sig0000007f : STD_LOGIC; 
  signal blk00000003_sig0000007e : STD_LOGIC; 
  signal blk00000003_sig0000007d : STD_LOGIC; 
  signal blk00000003_sig0000007c : STD_LOGIC; 
  signal blk00000003_sig0000007b : STD_LOGIC; 
  signal blk00000003_sig0000007a : STD_LOGIC; 
  signal blk00000003_sig00000079 : STD_LOGIC; 
  signal blk00000003_sig00000078 : STD_LOGIC; 
  signal blk00000003_sig00000077 : STD_LOGIC; 
  signal blk00000003_sig00000076 : STD_LOGIC; 
  signal blk00000003_sig00000075 : STD_LOGIC; 
  signal blk00000003_sig00000074 : STD_LOGIC; 
  signal blk00000003_sig00000073 : STD_LOGIC; 
  signal blk00000003_sig00000072 : STD_LOGIC; 
  signal blk00000003_sig00000071 : STD_LOGIC; 
  signal blk00000003_sig00000070 : STD_LOGIC; 
  signal blk00000003_sig0000006f : STD_LOGIC; 
  signal blk00000003_sig0000006e : STD_LOGIC; 
  signal blk00000003_sig0000006d : STD_LOGIC; 
  signal blk00000003_sig0000006c : STD_LOGIC; 
  signal blk00000003_sig0000006b : STD_LOGIC; 
  signal blk00000003_sig0000006a : STD_LOGIC; 
  signal blk00000003_sig00000069 : STD_LOGIC; 
  signal blk00000003_sig00000068 : STD_LOGIC; 
  signal blk00000003_sig00000067 : STD_LOGIC; 
  signal blk00000003_sig00000066 : STD_LOGIC; 
  signal blk00000003_sig00000065 : STD_LOGIC; 
  signal blk00000003_sig00000064 : STD_LOGIC; 
  signal blk00000003_sig00000063 : STD_LOGIC; 
  signal blk00000003_sig00000062 : STD_LOGIC; 
  signal blk00000003_sig00000061 : STD_LOGIC; 
  signal blk00000003_sig00000060 : STD_LOGIC; 
  signal blk00000003_sig0000005f : STD_LOGIC; 
  signal blk00000003_sig0000005e : STD_LOGIC; 
  signal blk00000003_sig0000005d : STD_LOGIC; 
  signal blk00000003_sig0000005c : STD_LOGIC; 
  signal blk00000003_sig0000005b : STD_LOGIC; 
  signal blk00000003_sig0000005a : STD_LOGIC; 
  signal blk00000003_sig00000059 : STD_LOGIC; 
  signal blk00000003_sig00000058 : STD_LOGIC; 
  signal blk00000003_sig00000057 : STD_LOGIC; 
  signal blk00000003_sig00000056 : STD_LOGIC; 
  signal blk00000003_sig00000055 : STD_LOGIC; 
  signal blk00000003_sig00000054 : STD_LOGIC; 
  signal blk00000003_sig00000053 : STD_LOGIC; 
  signal blk00000003_sig00000052 : STD_LOGIC; 
  signal blk00000003_sig00000051 : STD_LOGIC; 
  signal blk00000003_sig00000050 : STD_LOGIC; 
  signal blk00000003_sig0000004f : STD_LOGIC; 
  signal blk00000003_sig0000004e : STD_LOGIC; 
  signal blk00000003_sig0000004d : STD_LOGIC; 
  signal blk00000003_sig0000004c : STD_LOGIC; 
  signal blk00000003_sig0000004b : STD_LOGIC; 
  signal blk00000003_sig0000004a : STD_LOGIC; 
  signal blk00000003_sig00000049 : STD_LOGIC; 
  signal blk00000003_sig00000048 : STD_LOGIC; 
  signal blk00000003_sig00000047 : STD_LOGIC; 
  signal blk00000003_sig00000046 : STD_LOGIC; 
  signal blk00000003_sig00000045 : STD_LOGIC; 
  signal blk00000003_sig00000044 : STD_LOGIC; 
  signal blk00000003_sig00000043 : STD_LOGIC; 
  signal blk00000003_sig00000042 : STD_LOGIC; 
  signal blk00000003_sig00000041 : STD_LOGIC; 
  signal blk00000003_sig00000040 : STD_LOGIC; 
  signal blk00000003_sig0000003f : STD_LOGIC; 
  signal blk00000003_sig0000003e : STD_LOGIC; 
  signal blk00000003_sig0000003d : STD_LOGIC; 
  signal blk00000003_sig0000003c : STD_LOGIC; 
  signal blk00000003_sig0000003b : STD_LOGIC; 
  signal blk00000003_sig0000003a : STD_LOGIC; 
  signal blk00000003_sig00000039 : STD_LOGIC; 
  signal blk00000003_sig00000038 : STD_LOGIC; 
  signal blk00000003_sig00000037 : STD_LOGIC; 
  signal blk00000003_sig00000036 : STD_LOGIC; 
  signal blk00000003_sig00000035 : STD_LOGIC; 
  signal blk00000003_sig00000034 : STD_LOGIC; 
  signal blk00000003_sig00000033 : STD_LOGIC; 
  signal blk00000003_sig00000031 : STD_LOGIC; 
  signal NLW_blk00000001_P_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000002_G_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000003_blk0000032b_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000003_blk00000316_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000003_blk00000301_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000003_blk000002ec_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000003_blk000002d7_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000003_blk000002c2_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000003_blk000002ad_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000003_blk00000298_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000003_blk00000283_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000003_blk0000026e_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000003_blk00000259_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000003_blk00000244_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000003_blk0000022f_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000003_blk0000021a_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000003_blk00000205_O_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000003_blk000000fd_O_UNCONNECTED : STD_LOGIC; 
begin
  rfd <= NlwRenamedSig_OI_rfd;
  blk00000001 : VCC
    port map (
      P => NLW_blk00000001_P_UNCONNECTED
    );
  blk00000002 : GND
    port map (
      G => NLW_blk00000002_G_UNCONNECTED
    );
  blk00000003_blk000005e4 : INV
    port map (
      I => blk00000003_sig0000007e,
      O => blk00000003_sig00000130
    );
  blk00000003_blk000005e3 : INV
    port map (
      I => blk00000003_sig0000007d,
      O => blk00000003_sig00000133
    );
  blk00000003_blk000005e2 : INV
    port map (
      I => blk00000003_sig0000007c,
      O => blk00000003_sig00000136
    );
  blk00000003_blk000005e1 : INV
    port map (
      I => blk00000003_sig0000007b,
      O => blk00000003_sig00000139
    );
  blk00000003_blk000005e0 : INV
    port map (
      I => blk00000003_sig0000007a,
      O => blk00000003_sig0000013c
    );
  blk00000003_blk000005df : INV
    port map (
      I => blk00000003_sig000005ae,
      O => blk00000003_sig000005c9
    );
  blk00000003_blk000005de : INV
    port map (
      I => blk00000003_sig000005af,
      O => blk00000003_sig000005ca
    );
  blk00000003_blk000005dd : INV
    port map (
      I => blk00000003_sig000005b0,
      O => blk00000003_sig000005cb
    );
  blk00000003_blk000005dc : INV
    port map (
      I => blk00000003_sig000005b1,
      O => blk00000003_sig000005cc
    );
  blk00000003_blk000005db : INV
    port map (
      I => blk00000003_sig000005b2,
      O => blk00000003_sig000005cd
    );
  blk00000003_blk000005da : INV
    port map (
      I => blk00000003_sig000005b3,
      O => blk00000003_sig000005ce
    );
  blk00000003_blk000005d9 : INV
    port map (
      I => blk00000003_sig000005b4,
      O => blk00000003_sig000005cf
    );
  blk00000003_blk000005d8 : INV
    port map (
      I => blk00000003_sig000005b5,
      O => blk00000003_sig000005d0
    );
  blk00000003_blk000005d7 : INV
    port map (
      I => blk00000003_sig000005b6,
      O => blk00000003_sig000005d1
    );
  blk00000003_blk000005d6 : INV
    port map (
      I => blk00000003_sig000005b7,
      O => blk00000003_sig000005d2
    );
  blk00000003_blk000005d5 : INV
    port map (
      I => blk00000003_sig000005b8,
      O => blk00000003_sig000005d3
    );
  blk00000003_blk000005d4 : INV
    port map (
      I => blk00000003_sig000005b9,
      O => blk00000003_sig000005d4
    );
  blk00000003_blk000005d3 : INV
    port map (
      I => blk00000003_sig000005ba,
      O => blk00000003_sig000005d5
    );
  blk00000003_blk000005d2 : INV
    port map (
      I => blk00000003_sig000005bb,
      O => blk00000003_sig000005d6
    );
  blk00000003_blk000005d1 : INV
    port map (
      I => blk00000003_sig000005bc,
      O => blk00000003_sig000005d7
    );
  blk00000003_blk000005d0 : INV
    port map (
      I => blk00000003_sig000005bd,
      O => blk00000003_sig000005d8
    );
  blk00000003_blk000005cf : INV
    port map (
      I => blk00000003_sig000005be,
      O => blk00000003_sig000005d9
    );
  blk00000003_blk000005ce : INV
    port map (
      I => blk00000003_sig000005bf,
      O => blk00000003_sig000005da
    );
  blk00000003_blk000005cd : INV
    port map (
      I => blk00000003_sig000005c0,
      O => blk00000003_sig000005db
    );
  blk00000003_blk000005cc : INV
    port map (
      I => blk00000003_sig000005c1,
      O => blk00000003_sig000005dc
    );
  blk00000003_blk000005cb : INV
    port map (
      I => blk00000003_sig000005c2,
      O => blk00000003_sig000005dd
    );
  blk00000003_blk000005ca : INV
    port map (
      I => blk00000003_sig000005c3,
      O => blk00000003_sig000005de
    );
  blk00000003_blk000005c9 : INV
    port map (
      I => blk00000003_sig000005c4,
      O => blk00000003_sig000005df
    );
  blk00000003_blk000005c8 : INV
    port map (
      I => blk00000003_sig000005c5,
      O => blk00000003_sig000005e0
    );
  blk00000003_blk000005c7 : INV
    port map (
      I => blk00000003_sig000005c6,
      O => blk00000003_sig000005e1
    );
  blk00000003_blk000005c6 : INV
    port map (
      I => blk00000003_sig000005c7,
      O => blk00000003_sig000005e2
    );
  blk00000003_blk000005c5 : INV
    port map (
      I => blk00000003_sig000005c8,
      O => blk00000003_sig000005e3
    );
  blk00000003_blk000005c4 : INV
    port map (
      I => blk00000003_sig00000430,
      O => blk00000003_sig00000445
    );
  blk00000003_blk000005c3 : INV
    port map (
      I => blk00000003_sig00000414,
      O => blk00000003_sig00000429
    );
  blk00000003_blk000005c2 : INV
    port map (
      I => blk00000003_sig000003f8,
      O => blk00000003_sig0000040d
    );
  blk00000003_blk000005c1 : INV
    port map (
      I => blk00000003_sig000003dc,
      O => blk00000003_sig000003f1
    );
  blk00000003_blk000005c0 : INV
    port map (
      I => blk00000003_sig000003c0,
      O => blk00000003_sig000003d5
    );
  blk00000003_blk000005bf : INV
    port map (
      I => blk00000003_sig000003a4,
      O => blk00000003_sig000003b9
    );
  blk00000003_blk000005be : INV
    port map (
      I => blk00000003_sig00000388,
      O => blk00000003_sig0000039d
    );
  blk00000003_blk000005bd : INV
    port map (
      I => blk00000003_sig0000036c,
      O => blk00000003_sig00000381
    );
  blk00000003_blk000005bc : INV
    port map (
      I => blk00000003_sig00000350,
      O => blk00000003_sig00000365
    );
  blk00000003_blk000005bb : INV
    port map (
      I => blk00000003_sig00000334,
      O => blk00000003_sig00000349
    );
  blk00000003_blk000005ba : INV
    port map (
      I => blk00000003_sig00000318,
      O => blk00000003_sig0000032d
    );
  blk00000003_blk000005b9 : INV
    port map (
      I => blk00000003_sig000002fc,
      O => blk00000003_sig00000311
    );
  blk00000003_blk000005b8 : INV
    port map (
      I => blk00000003_sig000002e0,
      O => blk00000003_sig000002f5
    );
  blk00000003_blk000005b7 : INV
    port map (
      I => blk00000003_sig000002c4,
      O => blk00000003_sig000002d9
    );
  blk00000003_blk000005b6 : INV
    port map (
      I => blk00000003_sig000002a8,
      O => blk00000003_sig000002bd
    );
  blk00000003_blk000005b5 : INV
    port map (
      I => blk00000003_sig0000028c,
      O => blk00000003_sig000002a1
    );
  blk00000003_blk000005b4 : INV
    port map (
      I => blk00000003_sig0000026e,
      O => blk00000003_sig00000283
    );
  blk00000003_blk000005b3 : INV
    port map (
      I => blk00000003_sig00000250,
      O => blk00000003_sig00000265
    );
  blk00000003_blk000005b2 : INV
    port map (
      I => blk00000003_sig00000232,
      O => blk00000003_sig00000247
    );
  blk00000003_blk000005b1 : INV
    port map (
      I => blk00000003_sig00000214,
      O => blk00000003_sig00000229
    );
  blk00000003_blk000005b0 : INV
    port map (
      I => blk00000003_sig00000070,
      O => blk00000003_sig0000020b
    );
  blk00000003_blk000005af : INV
    port map (
      I => blk00000003_sig00000046,
      O => blk00000003_sig000001ee
    );
  blk00000003_blk000005ae : INV
    port map (
      I => blk00000003_sig00000059,
      O => blk00000003_sig000001d1
    );
  blk00000003_blk000005ad : INV
    port map (
      I => blk00000003_sig00000066,
      O => blk00000003_sig000001b3
    );
  blk00000003_blk000005ac : INV
    port map (
      I => blk00000003_sig0000006a,
      O => blk00000003_sig00000195
    );
  blk00000003_blk000005ab : INV
    port map (
      I => blk00000003_sig0000006d,
      O => blk00000003_sig00000177
    );
  blk00000003_blk000005aa : INV
    port map (
      I => blk00000003_sig0000006f,
      O => blk00000003_sig00000159
    );
  blk00000003_blk000005a9 : LUT1
    generic map(
      INIT => X"1"
    )
    port map (
      I0 => blk00000003_sig0000006f,
      O => blk00000003_sig000005e5
    );
  blk00000003_blk000005a8 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000042f,
      I1 => blk00000003_sig00000430,
      O => blk00000003_sig00000433
    );
  blk00000003_blk000005a7 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000042e,
      I1 => blk00000003_sig00000120,
      I2 => blk00000003_sig00000430,
      O => blk00000003_sig00000436
    );
  blk00000003_blk000005a6 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000042d,
      I1 => blk00000003_sig0000011f,
      I2 => blk00000003_sig00000430,
      O => blk00000003_sig00000439
    );
  blk00000003_blk000005a5 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000042c,
      I1 => blk00000003_sig0000011e,
      I2 => blk00000003_sig00000430,
      O => blk00000003_sig0000043c
    );
  blk00000003_blk000005a4 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000042b,
      I1 => blk00000003_sig0000011d,
      I2 => blk00000003_sig00000430,
      O => blk00000003_sig0000043f
    );
  blk00000003_blk000005a3 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000011b,
      I1 => blk00000003_sig0000011c,
      I2 => blk00000003_sig00000430,
      O => blk00000003_sig00000442
    );
  blk00000003_blk000005a2 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000011b,
      I1 => blk00000003_sig00000430,
      O => blk00000003_sig00000446
    );
  blk00000003_blk000005a1 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000413,
      I1 => blk00000003_sig00000414,
      O => blk00000003_sig00000417
    );
  blk00000003_blk000005a0 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000412,
      I1 => blk00000003_sig0000011a,
      I2 => blk00000003_sig00000414,
      O => blk00000003_sig0000041a
    );
  blk00000003_blk0000059f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000411,
      I1 => blk00000003_sig00000119,
      I2 => blk00000003_sig00000414,
      O => blk00000003_sig0000041d
    );
  blk00000003_blk0000059e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000410,
      I1 => blk00000003_sig00000118,
      I2 => blk00000003_sig00000414,
      O => blk00000003_sig00000420
    );
  blk00000003_blk0000059d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000040f,
      I1 => blk00000003_sig00000117,
      I2 => blk00000003_sig00000414,
      O => blk00000003_sig00000423
    );
  blk00000003_blk0000059c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000115,
      I1 => blk00000003_sig00000116,
      I2 => blk00000003_sig00000414,
      O => blk00000003_sig00000426
    );
  blk00000003_blk0000059b : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000115,
      I1 => blk00000003_sig00000414,
      O => blk00000003_sig0000042a
    );
  blk00000003_blk0000059a : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000003f7,
      I1 => blk00000003_sig000003f8,
      O => blk00000003_sig000003fb
    );
  blk00000003_blk00000599 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003f6,
      I1 => blk00000003_sig00000114,
      I2 => blk00000003_sig000003f8,
      O => blk00000003_sig000003fe
    );
  blk00000003_blk00000598 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003f5,
      I1 => blk00000003_sig00000113,
      I2 => blk00000003_sig000003f8,
      O => blk00000003_sig00000401
    );
  blk00000003_blk00000597 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003f4,
      I1 => blk00000003_sig00000112,
      I2 => blk00000003_sig000003f8,
      O => blk00000003_sig00000404
    );
  blk00000003_blk00000596 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003f3,
      I1 => blk00000003_sig00000111,
      I2 => blk00000003_sig000003f8,
      O => blk00000003_sig00000407
    );
  blk00000003_blk00000595 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000010f,
      I1 => blk00000003_sig00000110,
      I2 => blk00000003_sig000003f8,
      O => blk00000003_sig0000040a
    );
  blk00000003_blk00000594 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000010f,
      I1 => blk00000003_sig000003f8,
      O => blk00000003_sig0000040e
    );
  blk00000003_blk00000593 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000003db,
      I1 => blk00000003_sig000003dc,
      O => blk00000003_sig000003df
    );
  blk00000003_blk00000592 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003da,
      I1 => blk00000003_sig0000010e,
      I2 => blk00000003_sig000003dc,
      O => blk00000003_sig000003e2
    );
  blk00000003_blk00000591 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003d9,
      I1 => blk00000003_sig0000010d,
      I2 => blk00000003_sig000003dc,
      O => blk00000003_sig000003e5
    );
  blk00000003_blk00000590 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003d8,
      I1 => blk00000003_sig0000010c,
      I2 => blk00000003_sig000003dc,
      O => blk00000003_sig000003e8
    );
  blk00000003_blk0000058f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003d7,
      I1 => blk00000003_sig0000010b,
      I2 => blk00000003_sig000003dc,
      O => blk00000003_sig000003eb
    );
  blk00000003_blk0000058e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000109,
      I1 => blk00000003_sig0000010a,
      I2 => blk00000003_sig000003dc,
      O => blk00000003_sig000003ee
    );
  blk00000003_blk0000058d : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000109,
      I1 => blk00000003_sig000003dc,
      O => blk00000003_sig000003f2
    );
  blk00000003_blk0000058c : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000003bf,
      I1 => blk00000003_sig000003c0,
      O => blk00000003_sig000003c3
    );
  blk00000003_blk0000058b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003be,
      I1 => blk00000003_sig00000108,
      I2 => blk00000003_sig000003c0,
      O => blk00000003_sig000003c6
    );
  blk00000003_blk0000058a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003bd,
      I1 => blk00000003_sig00000107,
      I2 => blk00000003_sig000003c0,
      O => blk00000003_sig000003c9
    );
  blk00000003_blk00000589 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003bc,
      I1 => blk00000003_sig00000106,
      I2 => blk00000003_sig000003c0,
      O => blk00000003_sig000003cc
    );
  blk00000003_blk00000588 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003bb,
      I1 => blk00000003_sig00000105,
      I2 => blk00000003_sig000003c0,
      O => blk00000003_sig000003cf
    );
  blk00000003_blk00000587 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000103,
      I1 => blk00000003_sig00000104,
      I2 => blk00000003_sig000003c0,
      O => blk00000003_sig000003d2
    );
  blk00000003_blk00000586 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000103,
      I1 => blk00000003_sig000003c0,
      O => blk00000003_sig000003d6
    );
  blk00000003_blk00000585 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000003a3,
      I1 => blk00000003_sig000003a4,
      O => blk00000003_sig000003a7
    );
  blk00000003_blk00000584 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003a2,
      I1 => blk00000003_sig00000102,
      I2 => blk00000003_sig000003a4,
      O => blk00000003_sig000003aa
    );
  blk00000003_blk00000583 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003a1,
      I1 => blk00000003_sig00000101,
      I2 => blk00000003_sig000003a4,
      O => blk00000003_sig000003ad
    );
  blk00000003_blk00000582 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003a0,
      I1 => blk00000003_sig00000100,
      I2 => blk00000003_sig000003a4,
      O => blk00000003_sig000003b0
    );
  blk00000003_blk00000581 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000039f,
      I1 => blk00000003_sig000000ff,
      I2 => blk00000003_sig000003a4,
      O => blk00000003_sig000003b3
    );
  blk00000003_blk00000580 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000000fd,
      I1 => blk00000003_sig000000fe,
      I2 => blk00000003_sig000003a4,
      O => blk00000003_sig000003b6
    );
  blk00000003_blk0000057f : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000000fd,
      I1 => blk00000003_sig000003a4,
      O => blk00000003_sig000003ba
    );
  blk00000003_blk0000057e : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000387,
      I1 => blk00000003_sig00000388,
      O => blk00000003_sig0000038b
    );
  blk00000003_blk0000057d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000386,
      I1 => blk00000003_sig000000fc,
      I2 => blk00000003_sig00000388,
      O => blk00000003_sig0000038e
    );
  blk00000003_blk0000057c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000385,
      I1 => blk00000003_sig000000fb,
      I2 => blk00000003_sig00000388,
      O => blk00000003_sig00000391
    );
  blk00000003_blk0000057b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000384,
      I1 => blk00000003_sig000000fa,
      I2 => blk00000003_sig00000388,
      O => blk00000003_sig00000394
    );
  blk00000003_blk0000057a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000383,
      I1 => blk00000003_sig000000f9,
      I2 => blk00000003_sig00000388,
      O => blk00000003_sig00000397
    );
  blk00000003_blk00000579 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000000f7,
      I1 => blk00000003_sig000000f8,
      I2 => blk00000003_sig00000388,
      O => blk00000003_sig0000039a
    );
  blk00000003_blk00000578 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000000f7,
      I1 => blk00000003_sig00000388,
      O => blk00000003_sig0000039e
    );
  blk00000003_blk00000577 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000036b,
      I1 => blk00000003_sig0000036c,
      O => blk00000003_sig0000036f
    );
  blk00000003_blk00000576 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000036a,
      I1 => blk00000003_sig000000f6,
      I2 => blk00000003_sig0000036c,
      O => blk00000003_sig00000372
    );
  blk00000003_blk00000575 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000369,
      I1 => blk00000003_sig000000f5,
      I2 => blk00000003_sig0000036c,
      O => blk00000003_sig00000375
    );
  blk00000003_blk00000574 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000368,
      I1 => blk00000003_sig000000f4,
      I2 => blk00000003_sig0000036c,
      O => blk00000003_sig00000378
    );
  blk00000003_blk00000573 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000367,
      I1 => blk00000003_sig000000f3,
      I2 => blk00000003_sig0000036c,
      O => blk00000003_sig0000037b
    );
  blk00000003_blk00000572 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000000f1,
      I1 => blk00000003_sig000000f2,
      I2 => blk00000003_sig0000036c,
      O => blk00000003_sig0000037e
    );
  blk00000003_blk00000571 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000000f1,
      I1 => blk00000003_sig0000036c,
      O => blk00000003_sig00000382
    );
  blk00000003_blk00000570 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000034f,
      I1 => blk00000003_sig00000350,
      O => blk00000003_sig00000353
    );
  blk00000003_blk0000056f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000034e,
      I1 => blk00000003_sig000000f0,
      I2 => blk00000003_sig00000350,
      O => blk00000003_sig00000356
    );
  blk00000003_blk0000056e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000034d,
      I1 => blk00000003_sig000000ef,
      I2 => blk00000003_sig00000350,
      O => blk00000003_sig00000359
    );
  blk00000003_blk0000056d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000034c,
      I1 => blk00000003_sig000000ee,
      I2 => blk00000003_sig00000350,
      O => blk00000003_sig0000035c
    );
  blk00000003_blk0000056c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000034b,
      I1 => blk00000003_sig000000ed,
      I2 => blk00000003_sig00000350,
      O => blk00000003_sig0000035f
    );
  blk00000003_blk0000056b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000000eb,
      I1 => blk00000003_sig000000ec,
      I2 => blk00000003_sig00000350,
      O => blk00000003_sig00000362
    );
  blk00000003_blk0000056a : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000000eb,
      I1 => blk00000003_sig00000350,
      O => blk00000003_sig00000366
    );
  blk00000003_blk00000569 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000333,
      I1 => blk00000003_sig00000334,
      O => blk00000003_sig00000337
    );
  blk00000003_blk00000568 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000332,
      I1 => blk00000003_sig000000ea,
      I2 => blk00000003_sig00000334,
      O => blk00000003_sig0000033a
    );
  blk00000003_blk00000567 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000331,
      I1 => blk00000003_sig000000e9,
      I2 => blk00000003_sig00000334,
      O => blk00000003_sig0000033d
    );
  blk00000003_blk00000566 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000330,
      I1 => blk00000003_sig000000e8,
      I2 => blk00000003_sig00000334,
      O => blk00000003_sig00000340
    );
  blk00000003_blk00000565 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000032f,
      I1 => blk00000003_sig000000e7,
      I2 => blk00000003_sig00000334,
      O => blk00000003_sig00000343
    );
  blk00000003_blk00000564 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000000e5,
      I1 => blk00000003_sig000000e6,
      I2 => blk00000003_sig00000334,
      O => blk00000003_sig00000346
    );
  blk00000003_blk00000563 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000000e5,
      I1 => blk00000003_sig00000334,
      O => blk00000003_sig0000034a
    );
  blk00000003_blk00000562 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000317,
      I1 => blk00000003_sig00000318,
      O => blk00000003_sig0000031b
    );
  blk00000003_blk00000561 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000316,
      I1 => blk00000003_sig000000e4,
      I2 => blk00000003_sig00000318,
      O => blk00000003_sig0000031e
    );
  blk00000003_blk00000560 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000315,
      I1 => blk00000003_sig000000e3,
      I2 => blk00000003_sig00000318,
      O => blk00000003_sig00000321
    );
  blk00000003_blk0000055f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000314,
      I1 => blk00000003_sig000000e2,
      I2 => blk00000003_sig00000318,
      O => blk00000003_sig00000324
    );
  blk00000003_blk0000055e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000313,
      I1 => blk00000003_sig000000e1,
      I2 => blk00000003_sig00000318,
      O => blk00000003_sig00000327
    );
  blk00000003_blk0000055d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000000df,
      I1 => blk00000003_sig000000e0,
      I2 => blk00000003_sig00000318,
      O => blk00000003_sig0000032a
    );
  blk00000003_blk0000055c : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000000df,
      I1 => blk00000003_sig00000318,
      O => blk00000003_sig0000032e
    );
  blk00000003_blk0000055b : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000002fb,
      I1 => blk00000003_sig000002fc,
      O => blk00000003_sig000002ff
    );
  blk00000003_blk0000055a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002fa,
      I1 => blk00000003_sig000000de,
      I2 => blk00000003_sig000002fc,
      O => blk00000003_sig00000302
    );
  blk00000003_blk00000559 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002f9,
      I1 => blk00000003_sig000000dd,
      I2 => blk00000003_sig000002fc,
      O => blk00000003_sig00000305
    );
  blk00000003_blk00000558 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002f8,
      I1 => blk00000003_sig000000dc,
      I2 => blk00000003_sig000002fc,
      O => blk00000003_sig00000308
    );
  blk00000003_blk00000557 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002f7,
      I1 => blk00000003_sig000000db,
      I2 => blk00000003_sig000002fc,
      O => blk00000003_sig0000030b
    );
  blk00000003_blk00000556 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000000d9,
      I1 => blk00000003_sig000000da,
      I2 => blk00000003_sig000002fc,
      O => blk00000003_sig0000030e
    );
  blk00000003_blk00000555 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000000d9,
      I1 => blk00000003_sig000002fc,
      O => blk00000003_sig00000312
    );
  blk00000003_blk00000554 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000002df,
      I1 => blk00000003_sig000002e0,
      O => blk00000003_sig000002e3
    );
  blk00000003_blk00000553 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002de,
      I1 => blk00000003_sig000000d8,
      I2 => blk00000003_sig000002e0,
      O => blk00000003_sig000002e6
    );
  blk00000003_blk00000552 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002dd,
      I1 => blk00000003_sig000000d7,
      I2 => blk00000003_sig000002e0,
      O => blk00000003_sig000002e9
    );
  blk00000003_blk00000551 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002dc,
      I1 => blk00000003_sig000000d6,
      I2 => blk00000003_sig000002e0,
      O => blk00000003_sig000002ec
    );
  blk00000003_blk00000550 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002db,
      I1 => blk00000003_sig000000d5,
      I2 => blk00000003_sig000002e0,
      O => blk00000003_sig000002ef
    );
  blk00000003_blk0000054f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000000d3,
      I1 => blk00000003_sig000000d4,
      I2 => blk00000003_sig000002e0,
      O => blk00000003_sig000002f2
    );
  blk00000003_blk0000054e : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000000d3,
      I1 => blk00000003_sig000002e0,
      O => blk00000003_sig000002f6
    );
  blk00000003_blk0000054d : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000002c3,
      I1 => blk00000003_sig000002c4,
      O => blk00000003_sig000002c7
    );
  blk00000003_blk0000054c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002c2,
      I1 => blk00000003_sig000000d2,
      I2 => blk00000003_sig000002c4,
      O => blk00000003_sig000002ca
    );
  blk00000003_blk0000054b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002c1,
      I1 => blk00000003_sig000000d1,
      I2 => blk00000003_sig000002c4,
      O => blk00000003_sig000002cd
    );
  blk00000003_blk0000054a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002c0,
      I1 => blk00000003_sig000000d0,
      I2 => blk00000003_sig000002c4,
      O => blk00000003_sig000002d0
    );
  blk00000003_blk00000549 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002bf,
      I1 => blk00000003_sig000000cf,
      I2 => blk00000003_sig000002c4,
      O => blk00000003_sig000002d3
    );
  blk00000003_blk00000548 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000000cd,
      I1 => blk00000003_sig000000ce,
      I2 => blk00000003_sig000002c4,
      O => blk00000003_sig000002d6
    );
  blk00000003_blk00000547 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000000cd,
      I1 => blk00000003_sig000002c4,
      O => blk00000003_sig000002da
    );
  blk00000003_blk00000546 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000002a7,
      I1 => blk00000003_sig000002a8,
      O => blk00000003_sig000002ab
    );
  blk00000003_blk00000545 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002a6,
      I1 => blk00000003_sig000000cc,
      I2 => blk00000003_sig000002a8,
      O => blk00000003_sig000002ae
    );
  blk00000003_blk00000544 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002a5,
      I1 => blk00000003_sig000000cb,
      I2 => blk00000003_sig000002a8,
      O => blk00000003_sig000002b1
    );
  blk00000003_blk00000543 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002a4,
      I1 => blk00000003_sig000000ca,
      I2 => blk00000003_sig000002a8,
      O => blk00000003_sig000002b4
    );
  blk00000003_blk00000542 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002a3,
      I1 => blk00000003_sig000000c9,
      I2 => blk00000003_sig000002a8,
      O => blk00000003_sig000002b7
    );
  blk00000003_blk00000541 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000000c7,
      I1 => blk00000003_sig000000c8,
      I2 => blk00000003_sig000002a8,
      O => blk00000003_sig000002ba
    );
  blk00000003_blk00000540 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000000c7,
      I1 => blk00000003_sig000002a8,
      O => blk00000003_sig000002be
    );
  blk00000003_blk0000053f : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000028b,
      I1 => blk00000003_sig0000028c,
      O => blk00000003_sig0000028f
    );
  blk00000003_blk0000053e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000028a,
      I1 => blk00000003_sig000000c6,
      I2 => blk00000003_sig0000028c,
      O => blk00000003_sig00000292
    );
  blk00000003_blk0000053d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000289,
      I1 => blk00000003_sig000000c5,
      I2 => blk00000003_sig0000028c,
      O => blk00000003_sig00000295
    );
  blk00000003_blk0000053c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000288,
      I1 => blk00000003_sig000000c4,
      I2 => blk00000003_sig0000028c,
      O => blk00000003_sig00000298
    );
  blk00000003_blk0000053b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000287,
      I1 => blk00000003_sig000000c3,
      I2 => blk00000003_sig0000028c,
      O => blk00000003_sig0000029b
    );
  blk00000003_blk0000053a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000286,
      I1 => blk00000003_sig000000c2,
      I2 => blk00000003_sig0000028c,
      O => blk00000003_sig0000029e
    );
  blk00000003_blk00000539 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000000c1,
      I1 => blk00000003_sig0000028c,
      O => blk00000003_sig000002a2
    );
  blk00000003_blk00000538 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000026d,
      I1 => blk00000003_sig0000026e,
      O => blk00000003_sig00000271
    );
  blk00000003_blk00000537 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000026c,
      I1 => blk00000003_sig000000c0,
      I2 => blk00000003_sig0000026e,
      O => blk00000003_sig00000274
    );
  blk00000003_blk00000536 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000026b,
      I1 => blk00000003_sig000000bf,
      I2 => blk00000003_sig0000026e,
      O => blk00000003_sig00000277
    );
  blk00000003_blk00000535 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000026a,
      I1 => blk00000003_sig000000be,
      I2 => blk00000003_sig0000026e,
      O => blk00000003_sig0000027a
    );
  blk00000003_blk00000534 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000269,
      I1 => blk00000003_sig000000bd,
      I2 => blk00000003_sig0000026e,
      O => blk00000003_sig0000027d
    );
  blk00000003_blk00000533 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000268,
      I1 => blk00000003_sig000000bc,
      I2 => blk00000003_sig0000026e,
      O => blk00000003_sig00000280
    );
  blk00000003_blk00000532 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000078,
      I1 => blk00000003_sig000000bb,
      I2 => blk00000003_sig0000026e,
      O => blk00000003_sig00000284
    );
  blk00000003_blk00000531 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000024f,
      I1 => blk00000003_sig00000250,
      O => blk00000003_sig00000253
    );
  blk00000003_blk00000530 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000024e,
      I1 => blk00000003_sig000000ba,
      I2 => blk00000003_sig00000250,
      O => blk00000003_sig00000256
    );
  blk00000003_blk0000052f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000024d,
      I1 => blk00000003_sig000000b9,
      I2 => blk00000003_sig00000250,
      O => blk00000003_sig00000259
    );
  blk00000003_blk0000052e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000024c,
      I1 => blk00000003_sig000000b8,
      I2 => blk00000003_sig00000250,
      O => blk00000003_sig0000025c
    );
  blk00000003_blk0000052d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000024b,
      I1 => blk00000003_sig000000b7,
      I2 => blk00000003_sig00000250,
      O => blk00000003_sig0000025f
    );
  blk00000003_blk0000052c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000024a,
      I1 => blk00000003_sig000000b6,
      I2 => blk00000003_sig00000250,
      O => blk00000003_sig00000262
    );
  blk00000003_blk0000052b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000036,
      I1 => blk00000003_sig000000b5,
      I2 => blk00000003_sig00000250,
      O => blk00000003_sig00000266
    );
  blk00000003_blk0000052a : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000231,
      I1 => blk00000003_sig00000232,
      O => blk00000003_sig00000235
    );
  blk00000003_blk00000529 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000230,
      I1 => blk00000003_sig000000b4,
      I2 => blk00000003_sig00000232,
      O => blk00000003_sig00000238
    );
  blk00000003_blk00000528 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000022f,
      I1 => blk00000003_sig000000b3,
      I2 => blk00000003_sig00000232,
      O => blk00000003_sig0000023b
    );
  blk00000003_blk00000527 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000022e,
      I1 => blk00000003_sig000000b2,
      I2 => blk00000003_sig00000232,
      O => blk00000003_sig0000023e
    );
  blk00000003_blk00000526 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000022d,
      I1 => blk00000003_sig000000b1,
      I2 => blk00000003_sig00000232,
      O => blk00000003_sig00000241
    );
  blk00000003_blk00000525 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000022c,
      I1 => blk00000003_sig000000b0,
      I2 => blk00000003_sig00000232,
      O => blk00000003_sig00000244
    );
  blk00000003_blk00000524 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000003a,
      I1 => blk00000003_sig000000af,
      I2 => blk00000003_sig00000232,
      O => blk00000003_sig00000248
    );
  blk00000003_blk00000523 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000213,
      I1 => blk00000003_sig00000214,
      O => blk00000003_sig00000217
    );
  blk00000003_blk00000522 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000212,
      I1 => blk00000003_sig000000ae,
      I2 => blk00000003_sig00000214,
      O => blk00000003_sig0000021a
    );
  blk00000003_blk00000521 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000211,
      I1 => blk00000003_sig000000ad,
      I2 => blk00000003_sig00000214,
      O => blk00000003_sig0000021d
    );
  blk00000003_blk00000520 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000210,
      I1 => blk00000003_sig000000ac,
      I2 => blk00000003_sig00000214,
      O => blk00000003_sig00000220
    );
  blk00000003_blk0000051f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000020f,
      I1 => blk00000003_sig000000ab,
      I2 => blk00000003_sig00000214,
      O => blk00000003_sig00000223
    );
  blk00000003_blk0000051e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000020e,
      I1 => blk00000003_sig000000aa,
      I2 => blk00000003_sig00000214,
      O => blk00000003_sig00000226
    );
  blk00000003_blk0000051d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000003f,
      I1 => blk00000003_sig000000a9,
      I2 => blk00000003_sig00000214,
      O => blk00000003_sig0000022a
    );
  blk00000003_blk0000051c : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000001f6,
      I1 => blk00000003_sig00000070,
      O => blk00000003_sig000001f9
    );
  blk00000003_blk0000051b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001f5,
      I1 => blk00000003_sig000000a8,
      I2 => blk00000003_sig00000070,
      O => blk00000003_sig000001fc
    );
  blk00000003_blk0000051a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001f4,
      I1 => blk00000003_sig000000a7,
      I2 => blk00000003_sig00000070,
      O => blk00000003_sig000001ff
    );
  blk00000003_blk00000519 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001f3,
      I1 => blk00000003_sig000000a6,
      I2 => blk00000003_sig00000070,
      O => blk00000003_sig00000202
    );
  blk00000003_blk00000518 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001f2,
      I1 => blk00000003_sig000000a5,
      I2 => blk00000003_sig00000070,
      O => blk00000003_sig00000205
    );
  blk00000003_blk00000517 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001f1,
      I1 => blk00000003_sig000000a4,
      I2 => blk00000003_sig00000070,
      O => blk00000003_sig00000208
    );
  blk00000003_blk00000516 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000045,
      I1 => blk00000003_sig000000a3,
      I2 => blk00000003_sig00000070,
      O => blk00000003_sig0000020c
    );
  blk00000003_blk00000515 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000001d9,
      I1 => blk00000003_sig00000046,
      O => blk00000003_sig000001dc
    );
  blk00000003_blk00000514 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001d8,
      I1 => blk00000003_sig000000a2,
      I2 => blk00000003_sig00000046,
      O => blk00000003_sig000001df
    );
  blk00000003_blk00000513 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001d7,
      I1 => blk00000003_sig000000a1,
      I2 => blk00000003_sig00000046,
      O => blk00000003_sig000001e2
    );
  blk00000003_blk00000512 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001d6,
      I1 => blk00000003_sig000000a0,
      I2 => blk00000003_sig00000046,
      O => blk00000003_sig000001e5
    );
  blk00000003_blk00000511 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001d5,
      I1 => blk00000003_sig0000009f,
      I2 => blk00000003_sig00000046,
      O => blk00000003_sig000001e8
    );
  blk00000003_blk00000510 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001d4,
      I1 => blk00000003_sig0000009e,
      I2 => blk00000003_sig00000046,
      O => blk00000003_sig000001eb
    );
  blk00000003_blk0000050f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000058,
      I1 => blk00000003_sig0000009d,
      I2 => blk00000003_sig00000046,
      O => blk00000003_sig000001ef
    );
  blk00000003_blk0000050e : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000001bc,
      I1 => blk00000003_sig00000059,
      O => blk00000003_sig000001bf
    );
  blk00000003_blk0000050d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001bb,
      I1 => blk00000003_sig0000009c,
      I2 => blk00000003_sig00000059,
      O => blk00000003_sig000001c2
    );
  blk00000003_blk0000050c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001ba,
      I1 => blk00000003_sig0000009b,
      I2 => blk00000003_sig00000059,
      O => blk00000003_sig000001c5
    );
  blk00000003_blk0000050b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001b9,
      I1 => blk00000003_sig0000009a,
      I2 => blk00000003_sig00000059,
      O => blk00000003_sig000001c8
    );
  blk00000003_blk0000050a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001b8,
      I1 => blk00000003_sig00000099,
      I2 => blk00000003_sig00000059,
      O => blk00000003_sig000001cb
    );
  blk00000003_blk00000509 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001b7,
      I1 => blk00000003_sig00000098,
      I2 => blk00000003_sig00000059,
      O => blk00000003_sig000001ce
    );
  blk00000003_blk00000508 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000065,
      I1 => blk00000003_sig00000097,
      I2 => blk00000003_sig00000059,
      O => blk00000003_sig000001d2
    );
  blk00000003_blk00000507 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000019e,
      I1 => blk00000003_sig00000066,
      O => blk00000003_sig000001a1
    );
  blk00000003_blk00000506 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000019d,
      I1 => blk00000003_sig00000096,
      I2 => blk00000003_sig00000066,
      O => blk00000003_sig000001a4
    );
  blk00000003_blk00000505 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000019c,
      I1 => blk00000003_sig00000095,
      I2 => blk00000003_sig00000066,
      O => blk00000003_sig000001a7
    );
  blk00000003_blk00000504 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000019b,
      I1 => blk00000003_sig00000094,
      I2 => blk00000003_sig00000066,
      O => blk00000003_sig000001aa
    );
  blk00000003_blk00000503 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000019a,
      I1 => blk00000003_sig00000093,
      I2 => blk00000003_sig00000066,
      O => blk00000003_sig000001ad
    );
  blk00000003_blk00000502 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000199,
      I1 => blk00000003_sig00000092,
      I2 => blk00000003_sig00000066,
      O => blk00000003_sig000001b0
    );
  blk00000003_blk00000501 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001b6,
      I1 => blk00000003_sig00000091,
      I2 => blk00000003_sig00000066,
      O => blk00000003_sig000001b4
    );
  blk00000003_blk00000500 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000180,
      I1 => blk00000003_sig0000006a,
      O => blk00000003_sig00000183
    );
  blk00000003_blk000004ff : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000017f,
      I1 => blk00000003_sig00000090,
      I2 => blk00000003_sig0000006a,
      O => blk00000003_sig00000186
    );
  blk00000003_blk000004fe : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000017e,
      I1 => blk00000003_sig0000008f,
      I2 => blk00000003_sig0000006a,
      O => blk00000003_sig00000189
    );
  blk00000003_blk000004fd : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000017d,
      I1 => blk00000003_sig0000008e,
      I2 => blk00000003_sig0000006a,
      O => blk00000003_sig0000018c
    );
  blk00000003_blk000004fc : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000017c,
      I1 => blk00000003_sig0000008d,
      I2 => blk00000003_sig0000006a,
      O => blk00000003_sig0000018f
    );
  blk00000003_blk000004fb : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000017b,
      I1 => blk00000003_sig0000008c,
      I2 => blk00000003_sig0000006a,
      O => blk00000003_sig00000192
    );
  blk00000003_blk000004fa : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000198,
      I1 => blk00000003_sig0000008b,
      I2 => blk00000003_sig0000006a,
      O => blk00000003_sig00000196
    );
  blk00000003_blk000004f9 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000162,
      I1 => blk00000003_sig0000006d,
      O => blk00000003_sig00000165
    );
  blk00000003_blk000004f8 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000161,
      I1 => blk00000003_sig0000008a,
      I2 => blk00000003_sig0000006d,
      O => blk00000003_sig00000168
    );
  blk00000003_blk000004f7 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000160,
      I1 => blk00000003_sig00000089,
      I2 => blk00000003_sig0000006d,
      O => blk00000003_sig0000016b
    );
  blk00000003_blk000004f6 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000015f,
      I1 => blk00000003_sig00000088,
      I2 => blk00000003_sig0000006d,
      O => blk00000003_sig0000016e
    );
  blk00000003_blk000004f5 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000015e,
      I1 => blk00000003_sig00000087,
      I2 => blk00000003_sig0000006d,
      O => blk00000003_sig00000171
    );
  blk00000003_blk000004f4 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000015d,
      I1 => blk00000003_sig00000086,
      I2 => blk00000003_sig0000006d,
      O => blk00000003_sig00000174
    );
  blk00000003_blk000004f3 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000017a,
      I1 => blk00000003_sig00000085,
      I2 => blk00000003_sig0000006d,
      O => blk00000003_sig00000178
    );
  blk00000003_blk000004f2 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000145,
      I1 => blk00000003_sig0000006f,
      O => blk00000003_sig00000147
    );
  blk00000003_blk000004f1 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000144,
      I1 => blk00000003_sig00000084,
      I2 => blk00000003_sig0000006f,
      O => blk00000003_sig0000014a
    );
  blk00000003_blk000004f0 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000143,
      I1 => blk00000003_sig00000083,
      I2 => blk00000003_sig0000006f,
      O => blk00000003_sig0000014d
    );
  blk00000003_blk000004ef : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000142,
      I1 => blk00000003_sig00000082,
      I2 => blk00000003_sig0000006f,
      O => blk00000003_sig00000150
    );
  blk00000003_blk000004ee : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000141,
      I1 => blk00000003_sig00000081,
      I2 => blk00000003_sig0000006f,
      O => blk00000003_sig00000153
    );
  blk00000003_blk000004ed : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000140,
      I1 => blk00000003_sig00000080,
      I2 => blk00000003_sig0000006f,
      O => blk00000003_sig00000156
    );
  blk00000003_blk000004ec : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000015c,
      I1 => blk00000003_sig0000007f,
      I2 => blk00000003_sig0000006f,
      O => blk00000003_sig0000015a
    );
  blk00000003_blk000004eb : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000121,
      I1 => blk00000003_sig00000079,
      O => blk00000003_sig0000013e
    );
  blk00000003_blk000004ea : LUT1
    generic map(
      INIT => X"1"
    )
    port map (
      I0 => blk00000003_sig0000044e,
      O => blk00000003_sig000005e4
    );
  blk00000003_blk000004e9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005e4,
      Q => fractional(0)
    );
  blk00000003_blk000004e8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005e3,
      Q => fractional(1)
    );
  blk00000003_blk000004e7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005e2,
      Q => fractional(2)
    );
  blk00000003_blk000004e6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005e1,
      Q => fractional(3)
    );
  blk00000003_blk000004e5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005e0,
      Q => fractional(4)
    );
  blk00000003_blk000004e4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005df,
      Q => fractional(5)
    );
  blk00000003_blk000004e3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005de,
      Q => fractional(6)
    );
  blk00000003_blk000004e2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005dd,
      Q => fractional(7)
    );
  blk00000003_blk000004e1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005dc,
      Q => fractional(8)
    );
  blk00000003_blk000004e0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005db,
      Q => fractional(9)
    );
  blk00000003_blk000004df : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005da,
      Q => fractional(10)
    );
  blk00000003_blk000004de : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005d9,
      Q => fractional(11)
    );
  blk00000003_blk000004dd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005d8,
      Q => fractional(12)
    );
  blk00000003_blk000004dc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005d7,
      Q => fractional(13)
    );
  blk00000003_blk000004db : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005d6,
      Q => fractional(14)
    );
  blk00000003_blk000004da : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005d5,
      Q => fractional(15)
    );
  blk00000003_blk000004d9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005d4,
      Q => quotient(0)
    );
  blk00000003_blk000004d8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005d3,
      Q => quotient(1)
    );
  blk00000003_blk000004d7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005d2,
      Q => quotient(2)
    );
  blk00000003_blk000004d6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005d1,
      Q => quotient(3)
    );
  blk00000003_blk000004d5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005d0,
      Q => quotient(4)
    );
  blk00000003_blk000004d4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005cf,
      Q => quotient(5)
    );
  blk00000003_blk000004d3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005ce,
      Q => quotient(6)
    );
  blk00000003_blk000004d2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005cd,
      Q => quotient(7)
    );
  blk00000003_blk000004d1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005cc,
      Q => quotient(8)
    );
  blk00000003_blk000004d0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005cb,
      Q => quotient(9)
    );
  blk00000003_blk000004cf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005ca,
      Q => quotient(10)
    );
  blk00000003_blk000004ce : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005c9,
      Q => quotient(11)
    );
  blk00000003_blk000004cd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000430,
      Q => blk00000003_sig000005c8
    );
  blk00000003_blk000004cc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005ad,
      Q => blk00000003_sig000005c7
    );
  blk00000003_blk000004cb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005ac,
      Q => blk00000003_sig000005c6
    );
  blk00000003_blk000004ca : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005ab,
      Q => blk00000003_sig000005c5
    );
  blk00000003_blk000004c9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005aa,
      Q => blk00000003_sig000005c4
    );
  blk00000003_blk000004c8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005a9,
      Q => blk00000003_sig000005c3
    );
  blk00000003_blk000004c7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005a8,
      Q => blk00000003_sig000005c2
    );
  blk00000003_blk000004c6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005a7,
      Q => blk00000003_sig000005c1
    );
  blk00000003_blk000004c5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005a6,
      Q => blk00000003_sig000005c0
    );
  blk00000003_blk000004c4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005a5,
      Q => blk00000003_sig000005bf
    );
  blk00000003_blk000004c3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005a4,
      Q => blk00000003_sig000005be
    );
  blk00000003_blk000004c2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005a3,
      Q => blk00000003_sig000005bd
    );
  blk00000003_blk000004c1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005a2,
      Q => blk00000003_sig000005bc
    );
  blk00000003_blk000004c0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005a1,
      Q => blk00000003_sig000005bb
    );
  blk00000003_blk000004bf : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005a0,
      Q => blk00000003_sig000005ba
    );
  blk00000003_blk000004be : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000059f,
      Q => blk00000003_sig000005b9
    );
  blk00000003_blk000004bd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000059e,
      Q => blk00000003_sig000005b8
    );
  blk00000003_blk000004bc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000059d,
      Q => blk00000003_sig000005b7
    );
  blk00000003_blk000004bb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000059c,
      Q => blk00000003_sig000005b6
    );
  blk00000003_blk000004ba : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000059b,
      Q => blk00000003_sig000005b5
    );
  blk00000003_blk000004b9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000059a,
      Q => blk00000003_sig000005b4
    );
  blk00000003_blk000004b8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000599,
      Q => blk00000003_sig000005b3
    );
  blk00000003_blk000004b7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000598,
      Q => blk00000003_sig000005b2
    );
  blk00000003_blk000004b6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000597,
      Q => blk00000003_sig000005b1
    );
  blk00000003_blk000004b5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000596,
      Q => blk00000003_sig000005b0
    );
  blk00000003_blk000004b4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000595,
      Q => blk00000003_sig000005af
    );
  blk00000003_blk000004b3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000594,
      Q => blk00000003_sig000005ae
    );
  blk00000003_blk000004b2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000414,
      Q => blk00000003_sig000005ad
    );
  blk00000003_blk000004b1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000593,
      Q => blk00000003_sig000005ac
    );
  blk00000003_blk000004b0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000592,
      Q => blk00000003_sig000005ab
    );
  blk00000003_blk000004af : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000591,
      Q => blk00000003_sig000005aa
    );
  blk00000003_blk000004ae : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000590,
      Q => blk00000003_sig000005a9
    );
  blk00000003_blk000004ad : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000058f,
      Q => blk00000003_sig000005a8
    );
  blk00000003_blk000004ac : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000058e,
      Q => blk00000003_sig000005a7
    );
  blk00000003_blk000004ab : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000058d,
      Q => blk00000003_sig000005a6
    );
  blk00000003_blk000004aa : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000058c,
      Q => blk00000003_sig000005a5
    );
  blk00000003_blk000004a9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000058b,
      Q => blk00000003_sig000005a4
    );
  blk00000003_blk000004a8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000058a,
      Q => blk00000003_sig000005a3
    );
  blk00000003_blk000004a7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000589,
      Q => blk00000003_sig000005a2
    );
  blk00000003_blk000004a6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000588,
      Q => blk00000003_sig000005a1
    );
  blk00000003_blk000004a5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000587,
      Q => blk00000003_sig000005a0
    );
  blk00000003_blk000004a4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000586,
      Q => blk00000003_sig0000059f
    );
  blk00000003_blk000004a3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000585,
      Q => blk00000003_sig0000059e
    );
  blk00000003_blk000004a2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000584,
      Q => blk00000003_sig0000059d
    );
  blk00000003_blk000004a1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000583,
      Q => blk00000003_sig0000059c
    );
  blk00000003_blk000004a0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000582,
      Q => blk00000003_sig0000059b
    );
  blk00000003_blk0000049f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000581,
      Q => blk00000003_sig0000059a
    );
  blk00000003_blk0000049e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000580,
      Q => blk00000003_sig00000599
    );
  blk00000003_blk0000049d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000057f,
      Q => blk00000003_sig00000598
    );
  blk00000003_blk0000049c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000057e,
      Q => blk00000003_sig00000597
    );
  blk00000003_blk0000049b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000057d,
      Q => blk00000003_sig00000596
    );
  blk00000003_blk0000049a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000057c,
      Q => blk00000003_sig00000595
    );
  blk00000003_blk00000499 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000057b,
      Q => blk00000003_sig00000594
    );
  blk00000003_blk00000498 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003f8,
      Q => blk00000003_sig00000593
    );
  blk00000003_blk00000497 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000057a,
      Q => blk00000003_sig00000592
    );
  blk00000003_blk00000496 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000579,
      Q => blk00000003_sig00000591
    );
  blk00000003_blk00000495 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000578,
      Q => blk00000003_sig00000590
    );
  blk00000003_blk00000494 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000577,
      Q => blk00000003_sig0000058f
    );
  blk00000003_blk00000493 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000576,
      Q => blk00000003_sig0000058e
    );
  blk00000003_blk00000492 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000575,
      Q => blk00000003_sig0000058d
    );
  blk00000003_blk00000491 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000574,
      Q => blk00000003_sig0000058c
    );
  blk00000003_blk00000490 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000573,
      Q => blk00000003_sig0000058b
    );
  blk00000003_blk0000048f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000572,
      Q => blk00000003_sig0000058a
    );
  blk00000003_blk0000048e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000571,
      Q => blk00000003_sig00000589
    );
  blk00000003_blk0000048d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000570,
      Q => blk00000003_sig00000588
    );
  blk00000003_blk0000048c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000056f,
      Q => blk00000003_sig00000587
    );
  blk00000003_blk0000048b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000056e,
      Q => blk00000003_sig00000586
    );
  blk00000003_blk0000048a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000056d,
      Q => blk00000003_sig00000585
    );
  blk00000003_blk00000489 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000056c,
      Q => blk00000003_sig00000584
    );
  blk00000003_blk00000488 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000056b,
      Q => blk00000003_sig00000583
    );
  blk00000003_blk00000487 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000056a,
      Q => blk00000003_sig00000582
    );
  blk00000003_blk00000486 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000569,
      Q => blk00000003_sig00000581
    );
  blk00000003_blk00000485 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000568,
      Q => blk00000003_sig00000580
    );
  blk00000003_blk00000484 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000567,
      Q => blk00000003_sig0000057f
    );
  blk00000003_blk00000483 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000566,
      Q => blk00000003_sig0000057e
    );
  blk00000003_blk00000482 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000565,
      Q => blk00000003_sig0000057d
    );
  blk00000003_blk00000481 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000564,
      Q => blk00000003_sig0000057c
    );
  blk00000003_blk00000480 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000563,
      Q => blk00000003_sig0000057b
    );
  blk00000003_blk0000047f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003dc,
      Q => blk00000003_sig0000057a
    );
  blk00000003_blk0000047e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000562,
      Q => blk00000003_sig00000579
    );
  blk00000003_blk0000047d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000561,
      Q => blk00000003_sig00000578
    );
  blk00000003_blk0000047c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000560,
      Q => blk00000003_sig00000577
    );
  blk00000003_blk0000047b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000055f,
      Q => blk00000003_sig00000576
    );
  blk00000003_blk0000047a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000055e,
      Q => blk00000003_sig00000575
    );
  blk00000003_blk00000479 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000055d,
      Q => blk00000003_sig00000574
    );
  blk00000003_blk00000478 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000055c,
      Q => blk00000003_sig00000573
    );
  blk00000003_blk00000477 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000055b,
      Q => blk00000003_sig00000572
    );
  blk00000003_blk00000476 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000055a,
      Q => blk00000003_sig00000571
    );
  blk00000003_blk00000475 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000559,
      Q => blk00000003_sig00000570
    );
  blk00000003_blk00000474 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000558,
      Q => blk00000003_sig0000056f
    );
  blk00000003_blk00000473 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000557,
      Q => blk00000003_sig0000056e
    );
  blk00000003_blk00000472 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000556,
      Q => blk00000003_sig0000056d
    );
  blk00000003_blk00000471 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000555,
      Q => blk00000003_sig0000056c
    );
  blk00000003_blk00000470 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000554,
      Q => blk00000003_sig0000056b
    );
  blk00000003_blk0000046f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000553,
      Q => blk00000003_sig0000056a
    );
  blk00000003_blk0000046e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000552,
      Q => blk00000003_sig00000569
    );
  blk00000003_blk0000046d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000551,
      Q => blk00000003_sig00000568
    );
  blk00000003_blk0000046c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000550,
      Q => blk00000003_sig00000567
    );
  blk00000003_blk0000046b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000054f,
      Q => blk00000003_sig00000566
    );
  blk00000003_blk0000046a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000054e,
      Q => blk00000003_sig00000565
    );
  blk00000003_blk00000469 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000054d,
      Q => blk00000003_sig00000564
    );
  blk00000003_blk00000468 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000054c,
      Q => blk00000003_sig00000563
    );
  blk00000003_blk00000467 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003c0,
      Q => blk00000003_sig00000562
    );
  blk00000003_blk00000466 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000054b,
      Q => blk00000003_sig00000561
    );
  blk00000003_blk00000465 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000054a,
      Q => blk00000003_sig00000560
    );
  blk00000003_blk00000464 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000549,
      Q => blk00000003_sig0000055f
    );
  blk00000003_blk00000463 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000548,
      Q => blk00000003_sig0000055e
    );
  blk00000003_blk00000462 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000547,
      Q => blk00000003_sig0000055d
    );
  blk00000003_blk00000461 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000546,
      Q => blk00000003_sig0000055c
    );
  blk00000003_blk00000460 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000545,
      Q => blk00000003_sig0000055b
    );
  blk00000003_blk0000045f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000544,
      Q => blk00000003_sig0000055a
    );
  blk00000003_blk0000045e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000543,
      Q => blk00000003_sig00000559
    );
  blk00000003_blk0000045d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000542,
      Q => blk00000003_sig00000558
    );
  blk00000003_blk0000045c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000541,
      Q => blk00000003_sig00000557
    );
  blk00000003_blk0000045b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000540,
      Q => blk00000003_sig00000556
    );
  blk00000003_blk0000045a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000053f,
      Q => blk00000003_sig00000555
    );
  blk00000003_blk00000459 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000053e,
      Q => blk00000003_sig00000554
    );
  blk00000003_blk00000458 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000053d,
      Q => blk00000003_sig00000553
    );
  blk00000003_blk00000457 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000053c,
      Q => blk00000003_sig00000552
    );
  blk00000003_blk00000456 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000053b,
      Q => blk00000003_sig00000551
    );
  blk00000003_blk00000455 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000053a,
      Q => blk00000003_sig00000550
    );
  blk00000003_blk00000454 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000539,
      Q => blk00000003_sig0000054f
    );
  blk00000003_blk00000453 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000538,
      Q => blk00000003_sig0000054e
    );
  blk00000003_blk00000452 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000537,
      Q => blk00000003_sig0000054d
    );
  blk00000003_blk00000451 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000536,
      Q => blk00000003_sig0000054c
    );
  blk00000003_blk00000450 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003a4,
      Q => blk00000003_sig0000054b
    );
  blk00000003_blk0000044f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000535,
      Q => blk00000003_sig0000054a
    );
  blk00000003_blk0000044e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000534,
      Q => blk00000003_sig00000549
    );
  blk00000003_blk0000044d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000533,
      Q => blk00000003_sig00000548
    );
  blk00000003_blk0000044c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000532,
      Q => blk00000003_sig00000547
    );
  blk00000003_blk0000044b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000531,
      Q => blk00000003_sig00000546
    );
  blk00000003_blk0000044a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000530,
      Q => blk00000003_sig00000545
    );
  blk00000003_blk00000449 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000052f,
      Q => blk00000003_sig00000544
    );
  blk00000003_blk00000448 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000052e,
      Q => blk00000003_sig00000543
    );
  blk00000003_blk00000447 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000052d,
      Q => blk00000003_sig00000542
    );
  blk00000003_blk00000446 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000052c,
      Q => blk00000003_sig00000541
    );
  blk00000003_blk00000445 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000052b,
      Q => blk00000003_sig00000540
    );
  blk00000003_blk00000444 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000052a,
      Q => blk00000003_sig0000053f
    );
  blk00000003_blk00000443 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000529,
      Q => blk00000003_sig0000053e
    );
  blk00000003_blk00000442 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000528,
      Q => blk00000003_sig0000053d
    );
  blk00000003_blk00000441 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000527,
      Q => blk00000003_sig0000053c
    );
  blk00000003_blk00000440 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000526,
      Q => blk00000003_sig0000053b
    );
  blk00000003_blk0000043f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000525,
      Q => blk00000003_sig0000053a
    );
  blk00000003_blk0000043e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000524,
      Q => blk00000003_sig00000539
    );
  blk00000003_blk0000043d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000523,
      Q => blk00000003_sig00000538
    );
  blk00000003_blk0000043c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000522,
      Q => blk00000003_sig00000537
    );
  blk00000003_blk0000043b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000521,
      Q => blk00000003_sig00000536
    );
  blk00000003_blk0000043a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000388,
      Q => blk00000003_sig00000535
    );
  blk00000003_blk00000439 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000520,
      Q => blk00000003_sig00000534
    );
  blk00000003_blk00000438 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000051f,
      Q => blk00000003_sig00000533
    );
  blk00000003_blk00000437 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000051e,
      Q => blk00000003_sig00000532
    );
  blk00000003_blk00000436 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000051d,
      Q => blk00000003_sig00000531
    );
  blk00000003_blk00000435 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000051c,
      Q => blk00000003_sig00000530
    );
  blk00000003_blk00000434 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000051b,
      Q => blk00000003_sig0000052f
    );
  blk00000003_blk00000433 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000051a,
      Q => blk00000003_sig0000052e
    );
  blk00000003_blk00000432 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000519,
      Q => blk00000003_sig0000052d
    );
  blk00000003_blk00000431 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000518,
      Q => blk00000003_sig0000052c
    );
  blk00000003_blk00000430 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000517,
      Q => blk00000003_sig0000052b
    );
  blk00000003_blk0000042f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000516,
      Q => blk00000003_sig0000052a
    );
  blk00000003_blk0000042e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000515,
      Q => blk00000003_sig00000529
    );
  blk00000003_blk0000042d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000514,
      Q => blk00000003_sig00000528
    );
  blk00000003_blk0000042c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000513,
      Q => blk00000003_sig00000527
    );
  blk00000003_blk0000042b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000512,
      Q => blk00000003_sig00000526
    );
  blk00000003_blk0000042a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000511,
      Q => blk00000003_sig00000525
    );
  blk00000003_blk00000429 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000510,
      Q => blk00000003_sig00000524
    );
  blk00000003_blk00000428 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000050f,
      Q => blk00000003_sig00000523
    );
  blk00000003_blk00000427 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000050e,
      Q => blk00000003_sig00000522
    );
  blk00000003_blk00000426 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000050d,
      Q => blk00000003_sig00000521
    );
  blk00000003_blk00000425 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000036c,
      Q => blk00000003_sig00000520
    );
  blk00000003_blk00000424 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000050c,
      Q => blk00000003_sig0000051f
    );
  blk00000003_blk00000423 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000050b,
      Q => blk00000003_sig0000051e
    );
  blk00000003_blk00000422 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000050a,
      Q => blk00000003_sig0000051d
    );
  blk00000003_blk00000421 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000509,
      Q => blk00000003_sig0000051c
    );
  blk00000003_blk00000420 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000508,
      Q => blk00000003_sig0000051b
    );
  blk00000003_blk0000041f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000507,
      Q => blk00000003_sig0000051a
    );
  blk00000003_blk0000041e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000506,
      Q => blk00000003_sig00000519
    );
  blk00000003_blk0000041d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000505,
      Q => blk00000003_sig00000518
    );
  blk00000003_blk0000041c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000504,
      Q => blk00000003_sig00000517
    );
  blk00000003_blk0000041b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000503,
      Q => blk00000003_sig00000516
    );
  blk00000003_blk0000041a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000502,
      Q => blk00000003_sig00000515
    );
  blk00000003_blk00000419 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000501,
      Q => blk00000003_sig00000514
    );
  blk00000003_blk00000418 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000500,
      Q => blk00000003_sig00000513
    );
  blk00000003_blk00000417 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004ff,
      Q => blk00000003_sig00000512
    );
  blk00000003_blk00000416 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004fe,
      Q => blk00000003_sig00000511
    );
  blk00000003_blk00000415 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004fd,
      Q => blk00000003_sig00000510
    );
  blk00000003_blk00000414 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004fc,
      Q => blk00000003_sig0000050f
    );
  blk00000003_blk00000413 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004fb,
      Q => blk00000003_sig0000050e
    );
  blk00000003_blk00000412 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004fa,
      Q => blk00000003_sig0000050d
    );
  blk00000003_blk00000411 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000350,
      Q => blk00000003_sig0000050c
    );
  blk00000003_blk00000410 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004f9,
      Q => blk00000003_sig0000050b
    );
  blk00000003_blk0000040f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004f8,
      Q => blk00000003_sig0000050a
    );
  blk00000003_blk0000040e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004f7,
      Q => blk00000003_sig00000509
    );
  blk00000003_blk0000040d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004f6,
      Q => blk00000003_sig00000508
    );
  blk00000003_blk0000040c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004f5,
      Q => blk00000003_sig00000507
    );
  blk00000003_blk0000040b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004f4,
      Q => blk00000003_sig00000506
    );
  blk00000003_blk0000040a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004f3,
      Q => blk00000003_sig00000505
    );
  blk00000003_blk00000409 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004f2,
      Q => blk00000003_sig00000504
    );
  blk00000003_blk00000408 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004f1,
      Q => blk00000003_sig00000503
    );
  blk00000003_blk00000407 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004f0,
      Q => blk00000003_sig00000502
    );
  blk00000003_blk00000406 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004ef,
      Q => blk00000003_sig00000501
    );
  blk00000003_blk00000405 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004ee,
      Q => blk00000003_sig00000500
    );
  blk00000003_blk00000404 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004ed,
      Q => blk00000003_sig000004ff
    );
  blk00000003_blk00000403 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004ec,
      Q => blk00000003_sig000004fe
    );
  blk00000003_blk00000402 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004eb,
      Q => blk00000003_sig000004fd
    );
  blk00000003_blk00000401 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004ea,
      Q => blk00000003_sig000004fc
    );
  blk00000003_blk00000400 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004e9,
      Q => blk00000003_sig000004fb
    );
  blk00000003_blk000003ff : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004e8,
      Q => blk00000003_sig000004fa
    );
  blk00000003_blk000003fe : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000334,
      Q => blk00000003_sig000004f9
    );
  blk00000003_blk000003fd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004e7,
      Q => blk00000003_sig000004f8
    );
  blk00000003_blk000003fc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004e6,
      Q => blk00000003_sig000004f7
    );
  blk00000003_blk000003fb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004e5,
      Q => blk00000003_sig000004f6
    );
  blk00000003_blk000003fa : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004e4,
      Q => blk00000003_sig000004f5
    );
  blk00000003_blk000003f9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004e3,
      Q => blk00000003_sig000004f4
    );
  blk00000003_blk000003f8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004e2,
      Q => blk00000003_sig000004f3
    );
  blk00000003_blk000003f7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004e1,
      Q => blk00000003_sig000004f2
    );
  blk00000003_blk000003f6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004e0,
      Q => blk00000003_sig000004f1
    );
  blk00000003_blk000003f5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004df,
      Q => blk00000003_sig000004f0
    );
  blk00000003_blk000003f4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004de,
      Q => blk00000003_sig000004ef
    );
  blk00000003_blk000003f3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004dd,
      Q => blk00000003_sig000004ee
    );
  blk00000003_blk000003f2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004dc,
      Q => blk00000003_sig000004ed
    );
  blk00000003_blk000003f1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004db,
      Q => blk00000003_sig000004ec
    );
  blk00000003_blk000003f0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004da,
      Q => blk00000003_sig000004eb
    );
  blk00000003_blk000003ef : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004d9,
      Q => blk00000003_sig000004ea
    );
  blk00000003_blk000003ee : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004d8,
      Q => blk00000003_sig000004e9
    );
  blk00000003_blk000003ed : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004d7,
      Q => blk00000003_sig000004e8
    );
  blk00000003_blk000003ec : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000318,
      Q => blk00000003_sig000004e7
    );
  blk00000003_blk000003eb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004d6,
      Q => blk00000003_sig000004e6
    );
  blk00000003_blk000003ea : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004d5,
      Q => blk00000003_sig000004e5
    );
  blk00000003_blk000003e9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004d4,
      Q => blk00000003_sig000004e4
    );
  blk00000003_blk000003e8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004d3,
      Q => blk00000003_sig000004e3
    );
  blk00000003_blk000003e7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004d2,
      Q => blk00000003_sig000004e2
    );
  blk00000003_blk000003e6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004d1,
      Q => blk00000003_sig000004e1
    );
  blk00000003_blk000003e5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004d0,
      Q => blk00000003_sig000004e0
    );
  blk00000003_blk000003e4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004cf,
      Q => blk00000003_sig000004df
    );
  blk00000003_blk000003e3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004ce,
      Q => blk00000003_sig000004de
    );
  blk00000003_blk000003e2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004cd,
      Q => blk00000003_sig000004dd
    );
  blk00000003_blk000003e1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004cc,
      Q => blk00000003_sig000004dc
    );
  blk00000003_blk000003e0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004cb,
      Q => blk00000003_sig000004db
    );
  blk00000003_blk000003df : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004ca,
      Q => blk00000003_sig000004da
    );
  blk00000003_blk000003de : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004c9,
      Q => blk00000003_sig000004d9
    );
  blk00000003_blk000003dd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004c8,
      Q => blk00000003_sig000004d8
    );
  blk00000003_blk000003dc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004c7,
      Q => blk00000003_sig000004d7
    );
  blk00000003_blk000003db : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002fc,
      Q => blk00000003_sig000004d6
    );
  blk00000003_blk000003da : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004c6,
      Q => blk00000003_sig000004d5
    );
  blk00000003_blk000003d9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004c5,
      Q => blk00000003_sig000004d4
    );
  blk00000003_blk000003d8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004c4,
      Q => blk00000003_sig000004d3
    );
  blk00000003_blk000003d7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004c3,
      Q => blk00000003_sig000004d2
    );
  blk00000003_blk000003d6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004c2,
      Q => blk00000003_sig000004d1
    );
  blk00000003_blk000003d5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004c1,
      Q => blk00000003_sig000004d0
    );
  blk00000003_blk000003d4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004c0,
      Q => blk00000003_sig000004cf
    );
  blk00000003_blk000003d3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004bf,
      Q => blk00000003_sig000004ce
    );
  blk00000003_blk000003d2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004be,
      Q => blk00000003_sig000004cd
    );
  blk00000003_blk000003d1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004bd,
      Q => blk00000003_sig000004cc
    );
  blk00000003_blk000003d0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004bc,
      Q => blk00000003_sig000004cb
    );
  blk00000003_blk000003cf : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004bb,
      Q => blk00000003_sig000004ca
    );
  blk00000003_blk000003ce : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004ba,
      Q => blk00000003_sig000004c9
    );
  blk00000003_blk000003cd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004b9,
      Q => blk00000003_sig000004c8
    );
  blk00000003_blk000003cc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004b8,
      Q => blk00000003_sig000004c7
    );
  blk00000003_blk000003cb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002e0,
      Q => blk00000003_sig000004c6
    );
  blk00000003_blk000003ca : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004b7,
      Q => blk00000003_sig000004c5
    );
  blk00000003_blk000003c9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004b6,
      Q => blk00000003_sig000004c4
    );
  blk00000003_blk000003c8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004b5,
      Q => blk00000003_sig000004c3
    );
  blk00000003_blk000003c7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004b4,
      Q => blk00000003_sig000004c2
    );
  blk00000003_blk000003c6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004b3,
      Q => blk00000003_sig000004c1
    );
  blk00000003_blk000003c5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004b2,
      Q => blk00000003_sig000004c0
    );
  blk00000003_blk000003c4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004b1,
      Q => blk00000003_sig000004bf
    );
  blk00000003_blk000003c3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004b0,
      Q => blk00000003_sig000004be
    );
  blk00000003_blk000003c2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004af,
      Q => blk00000003_sig000004bd
    );
  blk00000003_blk000003c1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004ae,
      Q => blk00000003_sig000004bc
    );
  blk00000003_blk000003c0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004ad,
      Q => blk00000003_sig000004bb
    );
  blk00000003_blk000003bf : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004ac,
      Q => blk00000003_sig000004ba
    );
  blk00000003_blk000003be : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004ab,
      Q => blk00000003_sig000004b9
    );
  blk00000003_blk000003bd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004aa,
      Q => blk00000003_sig000004b8
    );
  blk00000003_blk000003bc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002c4,
      Q => blk00000003_sig000004b7
    );
  blk00000003_blk000003bb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004a9,
      Q => blk00000003_sig000004b6
    );
  blk00000003_blk000003ba : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004a8,
      Q => blk00000003_sig000004b5
    );
  blk00000003_blk000003b9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004a7,
      Q => blk00000003_sig000004b4
    );
  blk00000003_blk000003b8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004a6,
      Q => blk00000003_sig000004b3
    );
  blk00000003_blk000003b7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004a5,
      Q => blk00000003_sig000004b2
    );
  blk00000003_blk000003b6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004a4,
      Q => blk00000003_sig000004b1
    );
  blk00000003_blk000003b5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004a3,
      Q => blk00000003_sig000004b0
    );
  blk00000003_blk000003b4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004a2,
      Q => blk00000003_sig000004af
    );
  blk00000003_blk000003b3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004a1,
      Q => blk00000003_sig000004ae
    );
  blk00000003_blk000003b2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004a0,
      Q => blk00000003_sig000004ad
    );
  blk00000003_blk000003b1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000049f,
      Q => blk00000003_sig000004ac
    );
  blk00000003_blk000003b0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000049e,
      Q => blk00000003_sig000004ab
    );
  blk00000003_blk000003af : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000049d,
      Q => blk00000003_sig000004aa
    );
  blk00000003_blk000003ae : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002a8,
      Q => blk00000003_sig000004a9
    );
  blk00000003_blk000003ad : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000049c,
      Q => blk00000003_sig000004a8
    );
  blk00000003_blk000003ac : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000049b,
      Q => blk00000003_sig000004a7
    );
  blk00000003_blk000003ab : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000049a,
      Q => blk00000003_sig000004a6
    );
  blk00000003_blk000003aa : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000499,
      Q => blk00000003_sig000004a5
    );
  blk00000003_blk000003a9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000498,
      Q => blk00000003_sig000004a4
    );
  blk00000003_blk000003a8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000497,
      Q => blk00000003_sig000004a3
    );
  blk00000003_blk000003a7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000496,
      Q => blk00000003_sig000004a2
    );
  blk00000003_blk000003a6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000495,
      Q => blk00000003_sig000004a1
    );
  blk00000003_blk000003a5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000494,
      Q => blk00000003_sig000004a0
    );
  blk00000003_blk000003a4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000493,
      Q => blk00000003_sig0000049f
    );
  blk00000003_blk000003a3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000492,
      Q => blk00000003_sig0000049e
    );
  blk00000003_blk000003a2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000491,
      Q => blk00000003_sig0000049d
    );
  blk00000003_blk000003a1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000028c,
      Q => blk00000003_sig0000049c
    );
  blk00000003_blk000003a0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000490,
      Q => blk00000003_sig0000049b
    );
  blk00000003_blk0000039f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000048f,
      Q => blk00000003_sig0000049a
    );
  blk00000003_blk0000039e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000048e,
      Q => blk00000003_sig00000499
    );
  blk00000003_blk0000039d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000048d,
      Q => blk00000003_sig00000498
    );
  blk00000003_blk0000039c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000048c,
      Q => blk00000003_sig00000497
    );
  blk00000003_blk0000039b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000048b,
      Q => blk00000003_sig00000496
    );
  blk00000003_blk0000039a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000048a,
      Q => blk00000003_sig00000495
    );
  blk00000003_blk00000399 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000489,
      Q => blk00000003_sig00000494
    );
  blk00000003_blk00000398 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000488,
      Q => blk00000003_sig00000493
    );
  blk00000003_blk00000397 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000487,
      Q => blk00000003_sig00000492
    );
  blk00000003_blk00000396 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000486,
      Q => blk00000003_sig00000491
    );
  blk00000003_blk00000395 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000026e,
      Q => blk00000003_sig00000490
    );
  blk00000003_blk00000394 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000485,
      Q => blk00000003_sig0000048f
    );
  blk00000003_blk00000393 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000484,
      Q => blk00000003_sig0000048e
    );
  blk00000003_blk00000392 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000483,
      Q => blk00000003_sig0000048d
    );
  blk00000003_blk00000391 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000482,
      Q => blk00000003_sig0000048c
    );
  blk00000003_blk00000390 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000481,
      Q => blk00000003_sig0000048b
    );
  blk00000003_blk0000038f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000480,
      Q => blk00000003_sig0000048a
    );
  blk00000003_blk0000038e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000047f,
      Q => blk00000003_sig00000489
    );
  blk00000003_blk0000038d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000047e,
      Q => blk00000003_sig00000488
    );
  blk00000003_blk0000038c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000047d,
      Q => blk00000003_sig00000487
    );
  blk00000003_blk0000038b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000047c,
      Q => blk00000003_sig00000486
    );
  blk00000003_blk0000038a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000250,
      Q => blk00000003_sig00000485
    );
  blk00000003_blk00000389 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000047b,
      Q => blk00000003_sig00000484
    );
  blk00000003_blk00000388 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000047a,
      Q => blk00000003_sig00000483
    );
  blk00000003_blk00000387 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000479,
      Q => blk00000003_sig00000482
    );
  blk00000003_blk00000386 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000478,
      Q => blk00000003_sig00000481
    );
  blk00000003_blk00000385 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000477,
      Q => blk00000003_sig00000480
    );
  blk00000003_blk00000384 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000476,
      Q => blk00000003_sig0000047f
    );
  blk00000003_blk00000383 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000475,
      Q => blk00000003_sig0000047e
    );
  blk00000003_blk00000382 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000474,
      Q => blk00000003_sig0000047d
    );
  blk00000003_blk00000381 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000473,
      Q => blk00000003_sig0000047c
    );
  blk00000003_blk00000380 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000232,
      Q => blk00000003_sig0000047b
    );
  blk00000003_blk0000037f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000472,
      Q => blk00000003_sig0000047a
    );
  blk00000003_blk0000037e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000471,
      Q => blk00000003_sig00000479
    );
  blk00000003_blk0000037d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000470,
      Q => blk00000003_sig00000478
    );
  blk00000003_blk0000037c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000046f,
      Q => blk00000003_sig00000477
    );
  blk00000003_blk0000037b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000046e,
      Q => blk00000003_sig00000476
    );
  blk00000003_blk0000037a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000046d,
      Q => blk00000003_sig00000475
    );
  blk00000003_blk00000379 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000046c,
      Q => blk00000003_sig00000474
    );
  blk00000003_blk00000378 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000046b,
      Q => blk00000003_sig00000473
    );
  blk00000003_blk00000377 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000214,
      Q => blk00000003_sig00000472
    );
  blk00000003_blk00000376 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000071,
      Q => blk00000003_sig00000471
    );
  blk00000003_blk00000375 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000072,
      Q => blk00000003_sig00000470
    );
  blk00000003_blk00000374 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000073,
      Q => blk00000003_sig0000046f
    );
  blk00000003_blk00000373 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000074,
      Q => blk00000003_sig0000046e
    );
  blk00000003_blk00000372 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000075,
      Q => blk00000003_sig0000046d
    );
  blk00000003_blk00000371 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000076,
      Q => blk00000003_sig0000046c
    );
  blk00000003_blk00000370 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000077,
      Q => blk00000003_sig0000046b
    );
  blk00000003_blk0000036f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000046a,
      Q => blk00000003_sig0000005e
    );
  blk00000003_blk0000036e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000469,
      Q => blk00000003_sig0000005f
    );
  blk00000003_blk0000036d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000468,
      Q => blk00000003_sig00000060
    );
  blk00000003_blk0000036c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000467,
      Q => blk00000003_sig00000061
    );
  blk00000003_blk0000036b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000466,
      Q => blk00000003_sig00000062
    );
  blk00000003_blk0000036a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000465,
      Q => blk00000003_sig00000063
    );
  blk00000003_blk00000369 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000464,
      Q => blk00000003_sig00000064
    );
  blk00000003_blk00000368 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000463,
      Q => blk00000003_sig000001b6
    );
  blk00000003_blk00000367 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000462,
      Q => blk00000003_sig0000046a
    );
  blk00000003_blk00000366 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000461,
      Q => blk00000003_sig00000469
    );
  blk00000003_blk00000365 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000460,
      Q => blk00000003_sig00000468
    );
  blk00000003_blk00000364 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000045f,
      Q => blk00000003_sig00000467
    );
  blk00000003_blk00000363 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000045e,
      Q => blk00000003_sig00000466
    );
  blk00000003_blk00000362 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000045d,
      Q => blk00000003_sig00000465
    );
  blk00000003_blk00000361 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000045c,
      Q => blk00000003_sig00000464
    );
  blk00000003_blk00000360 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000045b,
      Q => blk00000003_sig00000463
    );
  blk00000003_blk0000035f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000045a,
      Q => blk00000003_sig00000198
    );
  blk00000003_blk0000035e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000459,
      Q => blk00000003_sig00000462
    );
  blk00000003_blk0000035d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000458,
      Q => blk00000003_sig00000461
    );
  blk00000003_blk0000035c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000457,
      Q => blk00000003_sig00000460
    );
  blk00000003_blk0000035b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000456,
      Q => blk00000003_sig0000045f
    );
  blk00000003_blk0000035a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000455,
      Q => blk00000003_sig0000045e
    );
  blk00000003_blk00000359 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000454,
      Q => blk00000003_sig0000045d
    );
  blk00000003_blk00000358 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000453,
      Q => blk00000003_sig0000045c
    );
  blk00000003_blk00000357 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000452,
      Q => blk00000003_sig0000045b
    );
  blk00000003_blk00000356 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000451,
      Q => blk00000003_sig0000045a
    );
  blk00000003_blk00000355 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000450,
      Q => blk00000003_sig0000017a
    );
  blk00000003_blk00000354 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000012c,
      Q => blk00000003_sig00000459
    );
  blk00000003_blk00000353 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000012b,
      Q => blk00000003_sig00000458
    );
  blk00000003_blk00000352 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000012a,
      Q => blk00000003_sig00000457
    );
  blk00000003_blk00000351 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000129,
      Q => blk00000003_sig00000456
    );
  blk00000003_blk00000350 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000128,
      Q => blk00000003_sig00000455
    );
  blk00000003_blk0000034f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000127,
      Q => blk00000003_sig00000454
    );
  blk00000003_blk0000034e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000126,
      Q => blk00000003_sig00000453
    );
  blk00000003_blk0000034d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000125,
      Q => blk00000003_sig00000452
    );
  blk00000003_blk0000034c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000124,
      Q => blk00000003_sig00000451
    );
  blk00000003_blk0000034b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000123,
      Q => blk00000003_sig00000450
    );
  blk00000003_blk0000034a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000122,
      Q => blk00000003_sig0000015c
    );
  blk00000003_blk00000349 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000444,
      Q => blk00000003_sig0000044f
    );
  blk00000003_blk00000348 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000434,
      Q => blk00000003_sig0000044e
    );
  blk00000003_blk00000347 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000437,
      Q => blk00000003_sig0000044d
    );
  blk00000003_blk00000346 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000043a,
      Q => blk00000003_sig0000044c
    );
  blk00000003_blk00000345 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000043d,
      Q => blk00000003_sig0000044b
    );
  blk00000003_blk00000344 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000440,
      Q => blk00000003_sig0000044a
    );
  blk00000003_blk00000343 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000443,
      Q => blk00000003_sig00000449
    );
  blk00000003_blk00000342 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000447,
      Q => blk00000003_sig00000448
    );
  blk00000003_blk00000341 : MUXCY
    port map (
      CI => blk00000003_sig00000445,
      DI => blk00000003_sig00000031,
      S => blk00000003_sig00000446,
      O => blk00000003_sig00000441
    );
  blk00000003_blk00000340 : XORCY
    port map (
      CI => blk00000003_sig00000445,
      LI => blk00000003_sig00000446,
      O => blk00000003_sig00000447
    );
  blk00000003_blk0000033f : MUXCY
    port map (
      CI => blk00000003_sig00000432,
      DI => blk00000003_sig0000042f,
      S => blk00000003_sig00000433,
      O => blk00000003_sig00000444
    );
  blk00000003_blk0000033e : MUXCY
    port map (
      CI => blk00000003_sig00000441,
      DI => blk00000003_sig0000011b,
      S => blk00000003_sig00000442,
      O => blk00000003_sig0000043e
    );
  blk00000003_blk0000033d : MUXCY
    port map (
      CI => blk00000003_sig0000043e,
      DI => blk00000003_sig0000042b,
      S => blk00000003_sig0000043f,
      O => blk00000003_sig0000043b
    );
  blk00000003_blk0000033c : MUXCY
    port map (
      CI => blk00000003_sig0000043b,
      DI => blk00000003_sig0000042c,
      S => blk00000003_sig0000043c,
      O => blk00000003_sig00000438
    );
  blk00000003_blk0000033b : MUXCY
    port map (
      CI => blk00000003_sig00000438,
      DI => blk00000003_sig0000042d,
      S => blk00000003_sig00000439,
      O => blk00000003_sig00000435
    );
  blk00000003_blk0000033a : MUXCY
    port map (
      CI => blk00000003_sig00000435,
      DI => blk00000003_sig0000042e,
      S => blk00000003_sig00000436,
      O => blk00000003_sig00000432
    );
  blk00000003_blk00000339 : XORCY
    port map (
      CI => blk00000003_sig00000441,
      LI => blk00000003_sig00000442,
      O => blk00000003_sig00000443
    );
  blk00000003_blk00000338 : XORCY
    port map (
      CI => blk00000003_sig0000043e,
      LI => blk00000003_sig0000043f,
      O => blk00000003_sig00000440
    );
  blk00000003_blk00000337 : XORCY
    port map (
      CI => blk00000003_sig0000043b,
      LI => blk00000003_sig0000043c,
      O => blk00000003_sig0000043d
    );
  blk00000003_blk00000336 : XORCY
    port map (
      CI => blk00000003_sig00000438,
      LI => blk00000003_sig00000439,
      O => blk00000003_sig0000043a
    );
  blk00000003_blk00000335 : XORCY
    port map (
      CI => blk00000003_sig00000435,
      LI => blk00000003_sig00000436,
      O => blk00000003_sig00000437
    );
  blk00000003_blk00000334 : XORCY
    port map (
      CI => blk00000003_sig00000432,
      LI => blk00000003_sig00000433,
      O => blk00000003_sig00000434
    );
  blk00000003_blk00000333 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000428,
      Q => blk00000003_sig00000431
    );
  blk00000003_blk00000332 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000418,
      Q => blk00000003_sig00000430
    );
  blk00000003_blk00000331 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000041b,
      Q => blk00000003_sig0000042f
    );
  blk00000003_blk00000330 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000041e,
      Q => blk00000003_sig0000042e
    );
  blk00000003_blk0000032f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000421,
      Q => blk00000003_sig0000042d
    );
  blk00000003_blk0000032e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000424,
      Q => blk00000003_sig0000042c
    );
  blk00000003_blk0000032d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000427,
      Q => blk00000003_sig0000042b
    );
  blk00000003_blk0000032c : MUXCY
    port map (
      CI => blk00000003_sig00000429,
      DI => blk00000003_sig00000031,
      S => blk00000003_sig0000042a,
      O => blk00000003_sig00000425
    );
  blk00000003_blk0000032b : XORCY
    port map (
      CI => blk00000003_sig00000429,
      LI => blk00000003_sig0000042a,
      O => NLW_blk00000003_blk0000032b_O_UNCONNECTED
    );
  blk00000003_blk0000032a : MUXCY
    port map (
      CI => blk00000003_sig00000416,
      DI => blk00000003_sig00000413,
      S => blk00000003_sig00000417,
      O => blk00000003_sig00000428
    );
  blk00000003_blk00000329 : MUXCY
    port map (
      CI => blk00000003_sig00000425,
      DI => blk00000003_sig00000115,
      S => blk00000003_sig00000426,
      O => blk00000003_sig00000422
    );
  blk00000003_blk00000328 : MUXCY
    port map (
      CI => blk00000003_sig00000422,
      DI => blk00000003_sig0000040f,
      S => blk00000003_sig00000423,
      O => blk00000003_sig0000041f
    );
  blk00000003_blk00000327 : MUXCY
    port map (
      CI => blk00000003_sig0000041f,
      DI => blk00000003_sig00000410,
      S => blk00000003_sig00000420,
      O => blk00000003_sig0000041c
    );
  blk00000003_blk00000326 : MUXCY
    port map (
      CI => blk00000003_sig0000041c,
      DI => blk00000003_sig00000411,
      S => blk00000003_sig0000041d,
      O => blk00000003_sig00000419
    );
  blk00000003_blk00000325 : MUXCY
    port map (
      CI => blk00000003_sig00000419,
      DI => blk00000003_sig00000412,
      S => blk00000003_sig0000041a,
      O => blk00000003_sig00000416
    );
  blk00000003_blk00000324 : XORCY
    port map (
      CI => blk00000003_sig00000425,
      LI => blk00000003_sig00000426,
      O => blk00000003_sig00000427
    );
  blk00000003_blk00000323 : XORCY
    port map (
      CI => blk00000003_sig00000422,
      LI => blk00000003_sig00000423,
      O => blk00000003_sig00000424
    );
  blk00000003_blk00000322 : XORCY
    port map (
      CI => blk00000003_sig0000041f,
      LI => blk00000003_sig00000420,
      O => blk00000003_sig00000421
    );
  blk00000003_blk00000321 : XORCY
    port map (
      CI => blk00000003_sig0000041c,
      LI => blk00000003_sig0000041d,
      O => blk00000003_sig0000041e
    );
  blk00000003_blk00000320 : XORCY
    port map (
      CI => blk00000003_sig00000419,
      LI => blk00000003_sig0000041a,
      O => blk00000003_sig0000041b
    );
  blk00000003_blk0000031f : XORCY
    port map (
      CI => blk00000003_sig00000416,
      LI => blk00000003_sig00000417,
      O => blk00000003_sig00000418
    );
  blk00000003_blk0000031e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000040c,
      Q => blk00000003_sig00000415
    );
  blk00000003_blk0000031d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003fc,
      Q => blk00000003_sig00000414
    );
  blk00000003_blk0000031c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003ff,
      Q => blk00000003_sig00000413
    );
  blk00000003_blk0000031b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000402,
      Q => blk00000003_sig00000412
    );
  blk00000003_blk0000031a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000405,
      Q => blk00000003_sig00000411
    );
  blk00000003_blk00000319 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000408,
      Q => blk00000003_sig00000410
    );
  blk00000003_blk00000318 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000040b,
      Q => blk00000003_sig0000040f
    );
  blk00000003_blk00000317 : MUXCY
    port map (
      CI => blk00000003_sig0000040d,
      DI => blk00000003_sig00000031,
      S => blk00000003_sig0000040e,
      O => blk00000003_sig00000409
    );
  blk00000003_blk00000316 : XORCY
    port map (
      CI => blk00000003_sig0000040d,
      LI => blk00000003_sig0000040e,
      O => NLW_blk00000003_blk00000316_O_UNCONNECTED
    );
  blk00000003_blk00000315 : MUXCY
    port map (
      CI => blk00000003_sig000003fa,
      DI => blk00000003_sig000003f7,
      S => blk00000003_sig000003fb,
      O => blk00000003_sig0000040c
    );
  blk00000003_blk00000314 : MUXCY
    port map (
      CI => blk00000003_sig00000409,
      DI => blk00000003_sig0000010f,
      S => blk00000003_sig0000040a,
      O => blk00000003_sig00000406
    );
  blk00000003_blk00000313 : MUXCY
    port map (
      CI => blk00000003_sig00000406,
      DI => blk00000003_sig000003f3,
      S => blk00000003_sig00000407,
      O => blk00000003_sig00000403
    );
  blk00000003_blk00000312 : MUXCY
    port map (
      CI => blk00000003_sig00000403,
      DI => blk00000003_sig000003f4,
      S => blk00000003_sig00000404,
      O => blk00000003_sig00000400
    );
  blk00000003_blk00000311 : MUXCY
    port map (
      CI => blk00000003_sig00000400,
      DI => blk00000003_sig000003f5,
      S => blk00000003_sig00000401,
      O => blk00000003_sig000003fd
    );
  blk00000003_blk00000310 : MUXCY
    port map (
      CI => blk00000003_sig000003fd,
      DI => blk00000003_sig000003f6,
      S => blk00000003_sig000003fe,
      O => blk00000003_sig000003fa
    );
  blk00000003_blk0000030f : XORCY
    port map (
      CI => blk00000003_sig00000409,
      LI => blk00000003_sig0000040a,
      O => blk00000003_sig0000040b
    );
  blk00000003_blk0000030e : XORCY
    port map (
      CI => blk00000003_sig00000406,
      LI => blk00000003_sig00000407,
      O => blk00000003_sig00000408
    );
  blk00000003_blk0000030d : XORCY
    port map (
      CI => blk00000003_sig00000403,
      LI => blk00000003_sig00000404,
      O => blk00000003_sig00000405
    );
  blk00000003_blk0000030c : XORCY
    port map (
      CI => blk00000003_sig00000400,
      LI => blk00000003_sig00000401,
      O => blk00000003_sig00000402
    );
  blk00000003_blk0000030b : XORCY
    port map (
      CI => blk00000003_sig000003fd,
      LI => blk00000003_sig000003fe,
      O => blk00000003_sig000003ff
    );
  blk00000003_blk0000030a : XORCY
    port map (
      CI => blk00000003_sig000003fa,
      LI => blk00000003_sig000003fb,
      O => blk00000003_sig000003fc
    );
  blk00000003_blk00000309 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003f0,
      Q => blk00000003_sig000003f9
    );
  blk00000003_blk00000308 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003e0,
      Q => blk00000003_sig000003f8
    );
  blk00000003_blk00000307 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003e3,
      Q => blk00000003_sig000003f7
    );
  blk00000003_blk00000306 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003e6,
      Q => blk00000003_sig000003f6
    );
  blk00000003_blk00000305 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003e9,
      Q => blk00000003_sig000003f5
    );
  blk00000003_blk00000304 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003ec,
      Q => blk00000003_sig000003f4
    );
  blk00000003_blk00000303 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003ef,
      Q => blk00000003_sig000003f3
    );
  blk00000003_blk00000302 : MUXCY
    port map (
      CI => blk00000003_sig000003f1,
      DI => blk00000003_sig00000031,
      S => blk00000003_sig000003f2,
      O => blk00000003_sig000003ed
    );
  blk00000003_blk00000301 : XORCY
    port map (
      CI => blk00000003_sig000003f1,
      LI => blk00000003_sig000003f2,
      O => NLW_blk00000003_blk00000301_O_UNCONNECTED
    );
  blk00000003_blk00000300 : MUXCY
    port map (
      CI => blk00000003_sig000003de,
      DI => blk00000003_sig000003db,
      S => blk00000003_sig000003df,
      O => blk00000003_sig000003f0
    );
  blk00000003_blk000002ff : MUXCY
    port map (
      CI => blk00000003_sig000003ed,
      DI => blk00000003_sig00000109,
      S => blk00000003_sig000003ee,
      O => blk00000003_sig000003ea
    );
  blk00000003_blk000002fe : MUXCY
    port map (
      CI => blk00000003_sig000003ea,
      DI => blk00000003_sig000003d7,
      S => blk00000003_sig000003eb,
      O => blk00000003_sig000003e7
    );
  blk00000003_blk000002fd : MUXCY
    port map (
      CI => blk00000003_sig000003e7,
      DI => blk00000003_sig000003d8,
      S => blk00000003_sig000003e8,
      O => blk00000003_sig000003e4
    );
  blk00000003_blk000002fc : MUXCY
    port map (
      CI => blk00000003_sig000003e4,
      DI => blk00000003_sig000003d9,
      S => blk00000003_sig000003e5,
      O => blk00000003_sig000003e1
    );
  blk00000003_blk000002fb : MUXCY
    port map (
      CI => blk00000003_sig000003e1,
      DI => blk00000003_sig000003da,
      S => blk00000003_sig000003e2,
      O => blk00000003_sig000003de
    );
  blk00000003_blk000002fa : XORCY
    port map (
      CI => blk00000003_sig000003ed,
      LI => blk00000003_sig000003ee,
      O => blk00000003_sig000003ef
    );
  blk00000003_blk000002f9 : XORCY
    port map (
      CI => blk00000003_sig000003ea,
      LI => blk00000003_sig000003eb,
      O => blk00000003_sig000003ec
    );
  blk00000003_blk000002f8 : XORCY
    port map (
      CI => blk00000003_sig000003e7,
      LI => blk00000003_sig000003e8,
      O => blk00000003_sig000003e9
    );
  blk00000003_blk000002f7 : XORCY
    port map (
      CI => blk00000003_sig000003e4,
      LI => blk00000003_sig000003e5,
      O => blk00000003_sig000003e6
    );
  blk00000003_blk000002f6 : XORCY
    port map (
      CI => blk00000003_sig000003e1,
      LI => blk00000003_sig000003e2,
      O => blk00000003_sig000003e3
    );
  blk00000003_blk000002f5 : XORCY
    port map (
      CI => blk00000003_sig000003de,
      LI => blk00000003_sig000003df,
      O => blk00000003_sig000003e0
    );
  blk00000003_blk000002f4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003d4,
      Q => blk00000003_sig000003dd
    );
  blk00000003_blk000002f3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003c4,
      Q => blk00000003_sig000003dc
    );
  blk00000003_blk000002f2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003c7,
      Q => blk00000003_sig000003db
    );
  blk00000003_blk000002f1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003ca,
      Q => blk00000003_sig000003da
    );
  blk00000003_blk000002f0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003cd,
      Q => blk00000003_sig000003d9
    );
  blk00000003_blk000002ef : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003d0,
      Q => blk00000003_sig000003d8
    );
  blk00000003_blk000002ee : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003d3,
      Q => blk00000003_sig000003d7
    );
  blk00000003_blk000002ed : MUXCY
    port map (
      CI => blk00000003_sig000003d5,
      DI => blk00000003_sig00000031,
      S => blk00000003_sig000003d6,
      O => blk00000003_sig000003d1
    );
  blk00000003_blk000002ec : XORCY
    port map (
      CI => blk00000003_sig000003d5,
      LI => blk00000003_sig000003d6,
      O => NLW_blk00000003_blk000002ec_O_UNCONNECTED
    );
  blk00000003_blk000002eb : MUXCY
    port map (
      CI => blk00000003_sig000003c2,
      DI => blk00000003_sig000003bf,
      S => blk00000003_sig000003c3,
      O => blk00000003_sig000003d4
    );
  blk00000003_blk000002ea : MUXCY
    port map (
      CI => blk00000003_sig000003d1,
      DI => blk00000003_sig00000103,
      S => blk00000003_sig000003d2,
      O => blk00000003_sig000003ce
    );
  blk00000003_blk000002e9 : MUXCY
    port map (
      CI => blk00000003_sig000003ce,
      DI => blk00000003_sig000003bb,
      S => blk00000003_sig000003cf,
      O => blk00000003_sig000003cb
    );
  blk00000003_blk000002e8 : MUXCY
    port map (
      CI => blk00000003_sig000003cb,
      DI => blk00000003_sig000003bc,
      S => blk00000003_sig000003cc,
      O => blk00000003_sig000003c8
    );
  blk00000003_blk000002e7 : MUXCY
    port map (
      CI => blk00000003_sig000003c8,
      DI => blk00000003_sig000003bd,
      S => blk00000003_sig000003c9,
      O => blk00000003_sig000003c5
    );
  blk00000003_blk000002e6 : MUXCY
    port map (
      CI => blk00000003_sig000003c5,
      DI => blk00000003_sig000003be,
      S => blk00000003_sig000003c6,
      O => blk00000003_sig000003c2
    );
  blk00000003_blk000002e5 : XORCY
    port map (
      CI => blk00000003_sig000003d1,
      LI => blk00000003_sig000003d2,
      O => blk00000003_sig000003d3
    );
  blk00000003_blk000002e4 : XORCY
    port map (
      CI => blk00000003_sig000003ce,
      LI => blk00000003_sig000003cf,
      O => blk00000003_sig000003d0
    );
  blk00000003_blk000002e3 : XORCY
    port map (
      CI => blk00000003_sig000003cb,
      LI => blk00000003_sig000003cc,
      O => blk00000003_sig000003cd
    );
  blk00000003_blk000002e2 : XORCY
    port map (
      CI => blk00000003_sig000003c8,
      LI => blk00000003_sig000003c9,
      O => blk00000003_sig000003ca
    );
  blk00000003_blk000002e1 : XORCY
    port map (
      CI => blk00000003_sig000003c5,
      LI => blk00000003_sig000003c6,
      O => blk00000003_sig000003c7
    );
  blk00000003_blk000002e0 : XORCY
    port map (
      CI => blk00000003_sig000003c2,
      LI => blk00000003_sig000003c3,
      O => blk00000003_sig000003c4
    );
  blk00000003_blk000002df : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003b8,
      Q => blk00000003_sig000003c1
    );
  blk00000003_blk000002de : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003a8,
      Q => blk00000003_sig000003c0
    );
  blk00000003_blk000002dd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003ab,
      Q => blk00000003_sig000003bf
    );
  blk00000003_blk000002dc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003ae,
      Q => blk00000003_sig000003be
    );
  blk00000003_blk000002db : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003b1,
      Q => blk00000003_sig000003bd
    );
  blk00000003_blk000002da : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003b4,
      Q => blk00000003_sig000003bc
    );
  blk00000003_blk000002d9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003b7,
      Q => blk00000003_sig000003bb
    );
  blk00000003_blk000002d8 : MUXCY
    port map (
      CI => blk00000003_sig000003b9,
      DI => blk00000003_sig00000031,
      S => blk00000003_sig000003ba,
      O => blk00000003_sig000003b5
    );
  blk00000003_blk000002d7 : XORCY
    port map (
      CI => blk00000003_sig000003b9,
      LI => blk00000003_sig000003ba,
      O => NLW_blk00000003_blk000002d7_O_UNCONNECTED
    );
  blk00000003_blk000002d6 : MUXCY
    port map (
      CI => blk00000003_sig000003a6,
      DI => blk00000003_sig000003a3,
      S => blk00000003_sig000003a7,
      O => blk00000003_sig000003b8
    );
  blk00000003_blk000002d5 : MUXCY
    port map (
      CI => blk00000003_sig000003b5,
      DI => blk00000003_sig000000fd,
      S => blk00000003_sig000003b6,
      O => blk00000003_sig000003b2
    );
  blk00000003_blk000002d4 : MUXCY
    port map (
      CI => blk00000003_sig000003b2,
      DI => blk00000003_sig0000039f,
      S => blk00000003_sig000003b3,
      O => blk00000003_sig000003af
    );
  blk00000003_blk000002d3 : MUXCY
    port map (
      CI => blk00000003_sig000003af,
      DI => blk00000003_sig000003a0,
      S => blk00000003_sig000003b0,
      O => blk00000003_sig000003ac
    );
  blk00000003_blk000002d2 : MUXCY
    port map (
      CI => blk00000003_sig000003ac,
      DI => blk00000003_sig000003a1,
      S => blk00000003_sig000003ad,
      O => blk00000003_sig000003a9
    );
  blk00000003_blk000002d1 : MUXCY
    port map (
      CI => blk00000003_sig000003a9,
      DI => blk00000003_sig000003a2,
      S => blk00000003_sig000003aa,
      O => blk00000003_sig000003a6
    );
  blk00000003_blk000002d0 : XORCY
    port map (
      CI => blk00000003_sig000003b5,
      LI => blk00000003_sig000003b6,
      O => blk00000003_sig000003b7
    );
  blk00000003_blk000002cf : XORCY
    port map (
      CI => blk00000003_sig000003b2,
      LI => blk00000003_sig000003b3,
      O => blk00000003_sig000003b4
    );
  blk00000003_blk000002ce : XORCY
    port map (
      CI => blk00000003_sig000003af,
      LI => blk00000003_sig000003b0,
      O => blk00000003_sig000003b1
    );
  blk00000003_blk000002cd : XORCY
    port map (
      CI => blk00000003_sig000003ac,
      LI => blk00000003_sig000003ad,
      O => blk00000003_sig000003ae
    );
  blk00000003_blk000002cc : XORCY
    port map (
      CI => blk00000003_sig000003a9,
      LI => blk00000003_sig000003aa,
      O => blk00000003_sig000003ab
    );
  blk00000003_blk000002cb : XORCY
    port map (
      CI => blk00000003_sig000003a6,
      LI => blk00000003_sig000003a7,
      O => blk00000003_sig000003a8
    );
  blk00000003_blk000002ca : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000039c,
      Q => blk00000003_sig000003a5
    );
  blk00000003_blk000002c9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000038c,
      Q => blk00000003_sig000003a4
    );
  blk00000003_blk000002c8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000038f,
      Q => blk00000003_sig000003a3
    );
  blk00000003_blk000002c7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000392,
      Q => blk00000003_sig000003a2
    );
  blk00000003_blk000002c6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000395,
      Q => blk00000003_sig000003a1
    );
  blk00000003_blk000002c5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000398,
      Q => blk00000003_sig000003a0
    );
  blk00000003_blk000002c4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000039b,
      Q => blk00000003_sig0000039f
    );
  blk00000003_blk000002c3 : MUXCY
    port map (
      CI => blk00000003_sig0000039d,
      DI => blk00000003_sig00000031,
      S => blk00000003_sig0000039e,
      O => blk00000003_sig00000399
    );
  blk00000003_blk000002c2 : XORCY
    port map (
      CI => blk00000003_sig0000039d,
      LI => blk00000003_sig0000039e,
      O => NLW_blk00000003_blk000002c2_O_UNCONNECTED
    );
  blk00000003_blk000002c1 : MUXCY
    port map (
      CI => blk00000003_sig0000038a,
      DI => blk00000003_sig00000387,
      S => blk00000003_sig0000038b,
      O => blk00000003_sig0000039c
    );
  blk00000003_blk000002c0 : MUXCY
    port map (
      CI => blk00000003_sig00000399,
      DI => blk00000003_sig000000f7,
      S => blk00000003_sig0000039a,
      O => blk00000003_sig00000396
    );
  blk00000003_blk000002bf : MUXCY
    port map (
      CI => blk00000003_sig00000396,
      DI => blk00000003_sig00000383,
      S => blk00000003_sig00000397,
      O => blk00000003_sig00000393
    );
  blk00000003_blk000002be : MUXCY
    port map (
      CI => blk00000003_sig00000393,
      DI => blk00000003_sig00000384,
      S => blk00000003_sig00000394,
      O => blk00000003_sig00000390
    );
  blk00000003_blk000002bd : MUXCY
    port map (
      CI => blk00000003_sig00000390,
      DI => blk00000003_sig00000385,
      S => blk00000003_sig00000391,
      O => blk00000003_sig0000038d
    );
  blk00000003_blk000002bc : MUXCY
    port map (
      CI => blk00000003_sig0000038d,
      DI => blk00000003_sig00000386,
      S => blk00000003_sig0000038e,
      O => blk00000003_sig0000038a
    );
  blk00000003_blk000002bb : XORCY
    port map (
      CI => blk00000003_sig00000399,
      LI => blk00000003_sig0000039a,
      O => blk00000003_sig0000039b
    );
  blk00000003_blk000002ba : XORCY
    port map (
      CI => blk00000003_sig00000396,
      LI => blk00000003_sig00000397,
      O => blk00000003_sig00000398
    );
  blk00000003_blk000002b9 : XORCY
    port map (
      CI => blk00000003_sig00000393,
      LI => blk00000003_sig00000394,
      O => blk00000003_sig00000395
    );
  blk00000003_blk000002b8 : XORCY
    port map (
      CI => blk00000003_sig00000390,
      LI => blk00000003_sig00000391,
      O => blk00000003_sig00000392
    );
  blk00000003_blk000002b7 : XORCY
    port map (
      CI => blk00000003_sig0000038d,
      LI => blk00000003_sig0000038e,
      O => blk00000003_sig0000038f
    );
  blk00000003_blk000002b6 : XORCY
    port map (
      CI => blk00000003_sig0000038a,
      LI => blk00000003_sig0000038b,
      O => blk00000003_sig0000038c
    );
  blk00000003_blk000002b5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000380,
      Q => blk00000003_sig00000389
    );
  blk00000003_blk000002b4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000370,
      Q => blk00000003_sig00000388
    );
  blk00000003_blk000002b3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000373,
      Q => blk00000003_sig00000387
    );
  blk00000003_blk000002b2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000376,
      Q => blk00000003_sig00000386
    );
  blk00000003_blk000002b1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000379,
      Q => blk00000003_sig00000385
    );
  blk00000003_blk000002b0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000037c,
      Q => blk00000003_sig00000384
    );
  blk00000003_blk000002af : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000037f,
      Q => blk00000003_sig00000383
    );
  blk00000003_blk000002ae : MUXCY
    port map (
      CI => blk00000003_sig00000381,
      DI => blk00000003_sig00000031,
      S => blk00000003_sig00000382,
      O => blk00000003_sig0000037d
    );
  blk00000003_blk000002ad : XORCY
    port map (
      CI => blk00000003_sig00000381,
      LI => blk00000003_sig00000382,
      O => NLW_blk00000003_blk000002ad_O_UNCONNECTED
    );
  blk00000003_blk000002ac : MUXCY
    port map (
      CI => blk00000003_sig0000036e,
      DI => blk00000003_sig0000036b,
      S => blk00000003_sig0000036f,
      O => blk00000003_sig00000380
    );
  blk00000003_blk000002ab : MUXCY
    port map (
      CI => blk00000003_sig0000037d,
      DI => blk00000003_sig000000f1,
      S => blk00000003_sig0000037e,
      O => blk00000003_sig0000037a
    );
  blk00000003_blk000002aa : MUXCY
    port map (
      CI => blk00000003_sig0000037a,
      DI => blk00000003_sig00000367,
      S => blk00000003_sig0000037b,
      O => blk00000003_sig00000377
    );
  blk00000003_blk000002a9 : MUXCY
    port map (
      CI => blk00000003_sig00000377,
      DI => blk00000003_sig00000368,
      S => blk00000003_sig00000378,
      O => blk00000003_sig00000374
    );
  blk00000003_blk000002a8 : MUXCY
    port map (
      CI => blk00000003_sig00000374,
      DI => blk00000003_sig00000369,
      S => blk00000003_sig00000375,
      O => blk00000003_sig00000371
    );
  blk00000003_blk000002a7 : MUXCY
    port map (
      CI => blk00000003_sig00000371,
      DI => blk00000003_sig0000036a,
      S => blk00000003_sig00000372,
      O => blk00000003_sig0000036e
    );
  blk00000003_blk000002a6 : XORCY
    port map (
      CI => blk00000003_sig0000037d,
      LI => blk00000003_sig0000037e,
      O => blk00000003_sig0000037f
    );
  blk00000003_blk000002a5 : XORCY
    port map (
      CI => blk00000003_sig0000037a,
      LI => blk00000003_sig0000037b,
      O => blk00000003_sig0000037c
    );
  blk00000003_blk000002a4 : XORCY
    port map (
      CI => blk00000003_sig00000377,
      LI => blk00000003_sig00000378,
      O => blk00000003_sig00000379
    );
  blk00000003_blk000002a3 : XORCY
    port map (
      CI => blk00000003_sig00000374,
      LI => blk00000003_sig00000375,
      O => blk00000003_sig00000376
    );
  blk00000003_blk000002a2 : XORCY
    port map (
      CI => blk00000003_sig00000371,
      LI => blk00000003_sig00000372,
      O => blk00000003_sig00000373
    );
  blk00000003_blk000002a1 : XORCY
    port map (
      CI => blk00000003_sig0000036e,
      LI => blk00000003_sig0000036f,
      O => blk00000003_sig00000370
    );
  blk00000003_blk000002a0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000364,
      Q => blk00000003_sig0000036d
    );
  blk00000003_blk0000029f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000354,
      Q => blk00000003_sig0000036c
    );
  blk00000003_blk0000029e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000357,
      Q => blk00000003_sig0000036b
    );
  blk00000003_blk0000029d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000035a,
      Q => blk00000003_sig0000036a
    );
  blk00000003_blk0000029c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000035d,
      Q => blk00000003_sig00000369
    );
  blk00000003_blk0000029b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000360,
      Q => blk00000003_sig00000368
    );
  blk00000003_blk0000029a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000363,
      Q => blk00000003_sig00000367
    );
  blk00000003_blk00000299 : MUXCY
    port map (
      CI => blk00000003_sig00000365,
      DI => blk00000003_sig00000031,
      S => blk00000003_sig00000366,
      O => blk00000003_sig00000361
    );
  blk00000003_blk00000298 : XORCY
    port map (
      CI => blk00000003_sig00000365,
      LI => blk00000003_sig00000366,
      O => NLW_blk00000003_blk00000298_O_UNCONNECTED
    );
  blk00000003_blk00000297 : MUXCY
    port map (
      CI => blk00000003_sig00000352,
      DI => blk00000003_sig0000034f,
      S => blk00000003_sig00000353,
      O => blk00000003_sig00000364
    );
  blk00000003_blk00000296 : MUXCY
    port map (
      CI => blk00000003_sig00000361,
      DI => blk00000003_sig000000eb,
      S => blk00000003_sig00000362,
      O => blk00000003_sig0000035e
    );
  blk00000003_blk00000295 : MUXCY
    port map (
      CI => blk00000003_sig0000035e,
      DI => blk00000003_sig0000034b,
      S => blk00000003_sig0000035f,
      O => blk00000003_sig0000035b
    );
  blk00000003_blk00000294 : MUXCY
    port map (
      CI => blk00000003_sig0000035b,
      DI => blk00000003_sig0000034c,
      S => blk00000003_sig0000035c,
      O => blk00000003_sig00000358
    );
  blk00000003_blk00000293 : MUXCY
    port map (
      CI => blk00000003_sig00000358,
      DI => blk00000003_sig0000034d,
      S => blk00000003_sig00000359,
      O => blk00000003_sig00000355
    );
  blk00000003_blk00000292 : MUXCY
    port map (
      CI => blk00000003_sig00000355,
      DI => blk00000003_sig0000034e,
      S => blk00000003_sig00000356,
      O => blk00000003_sig00000352
    );
  blk00000003_blk00000291 : XORCY
    port map (
      CI => blk00000003_sig00000361,
      LI => blk00000003_sig00000362,
      O => blk00000003_sig00000363
    );
  blk00000003_blk00000290 : XORCY
    port map (
      CI => blk00000003_sig0000035e,
      LI => blk00000003_sig0000035f,
      O => blk00000003_sig00000360
    );
  blk00000003_blk0000028f : XORCY
    port map (
      CI => blk00000003_sig0000035b,
      LI => blk00000003_sig0000035c,
      O => blk00000003_sig0000035d
    );
  blk00000003_blk0000028e : XORCY
    port map (
      CI => blk00000003_sig00000358,
      LI => blk00000003_sig00000359,
      O => blk00000003_sig0000035a
    );
  blk00000003_blk0000028d : XORCY
    port map (
      CI => blk00000003_sig00000355,
      LI => blk00000003_sig00000356,
      O => blk00000003_sig00000357
    );
  blk00000003_blk0000028c : XORCY
    port map (
      CI => blk00000003_sig00000352,
      LI => blk00000003_sig00000353,
      O => blk00000003_sig00000354
    );
  blk00000003_blk0000028b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000348,
      Q => blk00000003_sig00000351
    );
  blk00000003_blk0000028a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000338,
      Q => blk00000003_sig00000350
    );
  blk00000003_blk00000289 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000033b,
      Q => blk00000003_sig0000034f
    );
  blk00000003_blk00000288 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000033e,
      Q => blk00000003_sig0000034e
    );
  blk00000003_blk00000287 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000341,
      Q => blk00000003_sig0000034d
    );
  blk00000003_blk00000286 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000344,
      Q => blk00000003_sig0000034c
    );
  blk00000003_blk00000285 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000347,
      Q => blk00000003_sig0000034b
    );
  blk00000003_blk00000284 : MUXCY
    port map (
      CI => blk00000003_sig00000349,
      DI => blk00000003_sig00000031,
      S => blk00000003_sig0000034a,
      O => blk00000003_sig00000345
    );
  blk00000003_blk00000283 : XORCY
    port map (
      CI => blk00000003_sig00000349,
      LI => blk00000003_sig0000034a,
      O => NLW_blk00000003_blk00000283_O_UNCONNECTED
    );
  blk00000003_blk00000282 : MUXCY
    port map (
      CI => blk00000003_sig00000336,
      DI => blk00000003_sig00000333,
      S => blk00000003_sig00000337,
      O => blk00000003_sig00000348
    );
  blk00000003_blk00000281 : MUXCY
    port map (
      CI => blk00000003_sig00000345,
      DI => blk00000003_sig000000e5,
      S => blk00000003_sig00000346,
      O => blk00000003_sig00000342
    );
  blk00000003_blk00000280 : MUXCY
    port map (
      CI => blk00000003_sig00000342,
      DI => blk00000003_sig0000032f,
      S => blk00000003_sig00000343,
      O => blk00000003_sig0000033f
    );
  blk00000003_blk0000027f : MUXCY
    port map (
      CI => blk00000003_sig0000033f,
      DI => blk00000003_sig00000330,
      S => blk00000003_sig00000340,
      O => blk00000003_sig0000033c
    );
  blk00000003_blk0000027e : MUXCY
    port map (
      CI => blk00000003_sig0000033c,
      DI => blk00000003_sig00000331,
      S => blk00000003_sig0000033d,
      O => blk00000003_sig00000339
    );
  blk00000003_blk0000027d : MUXCY
    port map (
      CI => blk00000003_sig00000339,
      DI => blk00000003_sig00000332,
      S => blk00000003_sig0000033a,
      O => blk00000003_sig00000336
    );
  blk00000003_blk0000027c : XORCY
    port map (
      CI => blk00000003_sig00000345,
      LI => blk00000003_sig00000346,
      O => blk00000003_sig00000347
    );
  blk00000003_blk0000027b : XORCY
    port map (
      CI => blk00000003_sig00000342,
      LI => blk00000003_sig00000343,
      O => blk00000003_sig00000344
    );
  blk00000003_blk0000027a : XORCY
    port map (
      CI => blk00000003_sig0000033f,
      LI => blk00000003_sig00000340,
      O => blk00000003_sig00000341
    );
  blk00000003_blk00000279 : XORCY
    port map (
      CI => blk00000003_sig0000033c,
      LI => blk00000003_sig0000033d,
      O => blk00000003_sig0000033e
    );
  blk00000003_blk00000278 : XORCY
    port map (
      CI => blk00000003_sig00000339,
      LI => blk00000003_sig0000033a,
      O => blk00000003_sig0000033b
    );
  blk00000003_blk00000277 : XORCY
    port map (
      CI => blk00000003_sig00000336,
      LI => blk00000003_sig00000337,
      O => blk00000003_sig00000338
    );
  blk00000003_blk00000276 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000032c,
      Q => blk00000003_sig00000335
    );
  blk00000003_blk00000275 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000031c,
      Q => blk00000003_sig00000334
    );
  blk00000003_blk00000274 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000031f,
      Q => blk00000003_sig00000333
    );
  blk00000003_blk00000273 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000322,
      Q => blk00000003_sig00000332
    );
  blk00000003_blk00000272 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000325,
      Q => blk00000003_sig00000331
    );
  blk00000003_blk00000271 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000328,
      Q => blk00000003_sig00000330
    );
  blk00000003_blk00000270 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000032b,
      Q => blk00000003_sig0000032f
    );
  blk00000003_blk0000026f : MUXCY
    port map (
      CI => blk00000003_sig0000032d,
      DI => blk00000003_sig00000031,
      S => blk00000003_sig0000032e,
      O => blk00000003_sig00000329
    );
  blk00000003_blk0000026e : XORCY
    port map (
      CI => blk00000003_sig0000032d,
      LI => blk00000003_sig0000032e,
      O => NLW_blk00000003_blk0000026e_O_UNCONNECTED
    );
  blk00000003_blk0000026d : MUXCY
    port map (
      CI => blk00000003_sig0000031a,
      DI => blk00000003_sig00000317,
      S => blk00000003_sig0000031b,
      O => blk00000003_sig0000032c
    );
  blk00000003_blk0000026c : MUXCY
    port map (
      CI => blk00000003_sig00000329,
      DI => blk00000003_sig000000df,
      S => blk00000003_sig0000032a,
      O => blk00000003_sig00000326
    );
  blk00000003_blk0000026b : MUXCY
    port map (
      CI => blk00000003_sig00000326,
      DI => blk00000003_sig00000313,
      S => blk00000003_sig00000327,
      O => blk00000003_sig00000323
    );
  blk00000003_blk0000026a : MUXCY
    port map (
      CI => blk00000003_sig00000323,
      DI => blk00000003_sig00000314,
      S => blk00000003_sig00000324,
      O => blk00000003_sig00000320
    );
  blk00000003_blk00000269 : MUXCY
    port map (
      CI => blk00000003_sig00000320,
      DI => blk00000003_sig00000315,
      S => blk00000003_sig00000321,
      O => blk00000003_sig0000031d
    );
  blk00000003_blk00000268 : MUXCY
    port map (
      CI => blk00000003_sig0000031d,
      DI => blk00000003_sig00000316,
      S => blk00000003_sig0000031e,
      O => blk00000003_sig0000031a
    );
  blk00000003_blk00000267 : XORCY
    port map (
      CI => blk00000003_sig00000329,
      LI => blk00000003_sig0000032a,
      O => blk00000003_sig0000032b
    );
  blk00000003_blk00000266 : XORCY
    port map (
      CI => blk00000003_sig00000326,
      LI => blk00000003_sig00000327,
      O => blk00000003_sig00000328
    );
  blk00000003_blk00000265 : XORCY
    port map (
      CI => blk00000003_sig00000323,
      LI => blk00000003_sig00000324,
      O => blk00000003_sig00000325
    );
  blk00000003_blk00000264 : XORCY
    port map (
      CI => blk00000003_sig00000320,
      LI => blk00000003_sig00000321,
      O => blk00000003_sig00000322
    );
  blk00000003_blk00000263 : XORCY
    port map (
      CI => blk00000003_sig0000031d,
      LI => blk00000003_sig0000031e,
      O => blk00000003_sig0000031f
    );
  blk00000003_blk00000262 : XORCY
    port map (
      CI => blk00000003_sig0000031a,
      LI => blk00000003_sig0000031b,
      O => blk00000003_sig0000031c
    );
  blk00000003_blk00000261 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000310,
      Q => blk00000003_sig00000319
    );
  blk00000003_blk00000260 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000300,
      Q => blk00000003_sig00000318
    );
  blk00000003_blk0000025f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000303,
      Q => blk00000003_sig00000317
    );
  blk00000003_blk0000025e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000306,
      Q => blk00000003_sig00000316
    );
  blk00000003_blk0000025d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000309,
      Q => blk00000003_sig00000315
    );
  blk00000003_blk0000025c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000030c,
      Q => blk00000003_sig00000314
    );
  blk00000003_blk0000025b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000030f,
      Q => blk00000003_sig00000313
    );
  blk00000003_blk0000025a : MUXCY
    port map (
      CI => blk00000003_sig00000311,
      DI => blk00000003_sig00000031,
      S => blk00000003_sig00000312,
      O => blk00000003_sig0000030d
    );
  blk00000003_blk00000259 : XORCY
    port map (
      CI => blk00000003_sig00000311,
      LI => blk00000003_sig00000312,
      O => NLW_blk00000003_blk00000259_O_UNCONNECTED
    );
  blk00000003_blk00000258 : MUXCY
    port map (
      CI => blk00000003_sig000002fe,
      DI => blk00000003_sig000002fb,
      S => blk00000003_sig000002ff,
      O => blk00000003_sig00000310
    );
  blk00000003_blk00000257 : MUXCY
    port map (
      CI => blk00000003_sig0000030d,
      DI => blk00000003_sig000000d9,
      S => blk00000003_sig0000030e,
      O => blk00000003_sig0000030a
    );
  blk00000003_blk00000256 : MUXCY
    port map (
      CI => blk00000003_sig0000030a,
      DI => blk00000003_sig000002f7,
      S => blk00000003_sig0000030b,
      O => blk00000003_sig00000307
    );
  blk00000003_blk00000255 : MUXCY
    port map (
      CI => blk00000003_sig00000307,
      DI => blk00000003_sig000002f8,
      S => blk00000003_sig00000308,
      O => blk00000003_sig00000304
    );
  blk00000003_blk00000254 : MUXCY
    port map (
      CI => blk00000003_sig00000304,
      DI => blk00000003_sig000002f9,
      S => blk00000003_sig00000305,
      O => blk00000003_sig00000301
    );
  blk00000003_blk00000253 : MUXCY
    port map (
      CI => blk00000003_sig00000301,
      DI => blk00000003_sig000002fa,
      S => blk00000003_sig00000302,
      O => blk00000003_sig000002fe
    );
  blk00000003_blk00000252 : XORCY
    port map (
      CI => blk00000003_sig0000030d,
      LI => blk00000003_sig0000030e,
      O => blk00000003_sig0000030f
    );
  blk00000003_blk00000251 : XORCY
    port map (
      CI => blk00000003_sig0000030a,
      LI => blk00000003_sig0000030b,
      O => blk00000003_sig0000030c
    );
  blk00000003_blk00000250 : XORCY
    port map (
      CI => blk00000003_sig00000307,
      LI => blk00000003_sig00000308,
      O => blk00000003_sig00000309
    );
  blk00000003_blk0000024f : XORCY
    port map (
      CI => blk00000003_sig00000304,
      LI => blk00000003_sig00000305,
      O => blk00000003_sig00000306
    );
  blk00000003_blk0000024e : XORCY
    port map (
      CI => blk00000003_sig00000301,
      LI => blk00000003_sig00000302,
      O => blk00000003_sig00000303
    );
  blk00000003_blk0000024d : XORCY
    port map (
      CI => blk00000003_sig000002fe,
      LI => blk00000003_sig000002ff,
      O => blk00000003_sig00000300
    );
  blk00000003_blk0000024c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002f4,
      Q => blk00000003_sig000002fd
    );
  blk00000003_blk0000024b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002e4,
      Q => blk00000003_sig000002fc
    );
  blk00000003_blk0000024a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002e7,
      Q => blk00000003_sig000002fb
    );
  blk00000003_blk00000249 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002ea,
      Q => blk00000003_sig000002fa
    );
  blk00000003_blk00000248 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002ed,
      Q => blk00000003_sig000002f9
    );
  blk00000003_blk00000247 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002f0,
      Q => blk00000003_sig000002f8
    );
  blk00000003_blk00000246 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002f3,
      Q => blk00000003_sig000002f7
    );
  blk00000003_blk00000245 : MUXCY
    port map (
      CI => blk00000003_sig000002f5,
      DI => blk00000003_sig00000031,
      S => blk00000003_sig000002f6,
      O => blk00000003_sig000002f1
    );
  blk00000003_blk00000244 : XORCY
    port map (
      CI => blk00000003_sig000002f5,
      LI => blk00000003_sig000002f6,
      O => NLW_blk00000003_blk00000244_O_UNCONNECTED
    );
  blk00000003_blk00000243 : MUXCY
    port map (
      CI => blk00000003_sig000002e2,
      DI => blk00000003_sig000002df,
      S => blk00000003_sig000002e3,
      O => blk00000003_sig000002f4
    );
  blk00000003_blk00000242 : MUXCY
    port map (
      CI => blk00000003_sig000002f1,
      DI => blk00000003_sig000000d3,
      S => blk00000003_sig000002f2,
      O => blk00000003_sig000002ee
    );
  blk00000003_blk00000241 : MUXCY
    port map (
      CI => blk00000003_sig000002ee,
      DI => blk00000003_sig000002db,
      S => blk00000003_sig000002ef,
      O => blk00000003_sig000002eb
    );
  blk00000003_blk00000240 : MUXCY
    port map (
      CI => blk00000003_sig000002eb,
      DI => blk00000003_sig000002dc,
      S => blk00000003_sig000002ec,
      O => blk00000003_sig000002e8
    );
  blk00000003_blk0000023f : MUXCY
    port map (
      CI => blk00000003_sig000002e8,
      DI => blk00000003_sig000002dd,
      S => blk00000003_sig000002e9,
      O => blk00000003_sig000002e5
    );
  blk00000003_blk0000023e : MUXCY
    port map (
      CI => blk00000003_sig000002e5,
      DI => blk00000003_sig000002de,
      S => blk00000003_sig000002e6,
      O => blk00000003_sig000002e2
    );
  blk00000003_blk0000023d : XORCY
    port map (
      CI => blk00000003_sig000002f1,
      LI => blk00000003_sig000002f2,
      O => blk00000003_sig000002f3
    );
  blk00000003_blk0000023c : XORCY
    port map (
      CI => blk00000003_sig000002ee,
      LI => blk00000003_sig000002ef,
      O => blk00000003_sig000002f0
    );
  blk00000003_blk0000023b : XORCY
    port map (
      CI => blk00000003_sig000002eb,
      LI => blk00000003_sig000002ec,
      O => blk00000003_sig000002ed
    );
  blk00000003_blk0000023a : XORCY
    port map (
      CI => blk00000003_sig000002e8,
      LI => blk00000003_sig000002e9,
      O => blk00000003_sig000002ea
    );
  blk00000003_blk00000239 : XORCY
    port map (
      CI => blk00000003_sig000002e5,
      LI => blk00000003_sig000002e6,
      O => blk00000003_sig000002e7
    );
  blk00000003_blk00000238 : XORCY
    port map (
      CI => blk00000003_sig000002e2,
      LI => blk00000003_sig000002e3,
      O => blk00000003_sig000002e4
    );
  blk00000003_blk00000237 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002d8,
      Q => blk00000003_sig000002e1
    );
  blk00000003_blk00000236 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002c8,
      Q => blk00000003_sig000002e0
    );
  blk00000003_blk00000235 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002cb,
      Q => blk00000003_sig000002df
    );
  blk00000003_blk00000234 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002ce,
      Q => blk00000003_sig000002de
    );
  blk00000003_blk00000233 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002d1,
      Q => blk00000003_sig000002dd
    );
  blk00000003_blk00000232 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002d4,
      Q => blk00000003_sig000002dc
    );
  blk00000003_blk00000231 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002d7,
      Q => blk00000003_sig000002db
    );
  blk00000003_blk00000230 : MUXCY
    port map (
      CI => blk00000003_sig000002d9,
      DI => blk00000003_sig00000031,
      S => blk00000003_sig000002da,
      O => blk00000003_sig000002d5
    );
  blk00000003_blk0000022f : XORCY
    port map (
      CI => blk00000003_sig000002d9,
      LI => blk00000003_sig000002da,
      O => NLW_blk00000003_blk0000022f_O_UNCONNECTED
    );
  blk00000003_blk0000022e : MUXCY
    port map (
      CI => blk00000003_sig000002c6,
      DI => blk00000003_sig000002c3,
      S => blk00000003_sig000002c7,
      O => blk00000003_sig000002d8
    );
  blk00000003_blk0000022d : MUXCY
    port map (
      CI => blk00000003_sig000002d5,
      DI => blk00000003_sig000000cd,
      S => blk00000003_sig000002d6,
      O => blk00000003_sig000002d2
    );
  blk00000003_blk0000022c : MUXCY
    port map (
      CI => blk00000003_sig000002d2,
      DI => blk00000003_sig000002bf,
      S => blk00000003_sig000002d3,
      O => blk00000003_sig000002cf
    );
  blk00000003_blk0000022b : MUXCY
    port map (
      CI => blk00000003_sig000002cf,
      DI => blk00000003_sig000002c0,
      S => blk00000003_sig000002d0,
      O => blk00000003_sig000002cc
    );
  blk00000003_blk0000022a : MUXCY
    port map (
      CI => blk00000003_sig000002cc,
      DI => blk00000003_sig000002c1,
      S => blk00000003_sig000002cd,
      O => blk00000003_sig000002c9
    );
  blk00000003_blk00000229 : MUXCY
    port map (
      CI => blk00000003_sig000002c9,
      DI => blk00000003_sig000002c2,
      S => blk00000003_sig000002ca,
      O => blk00000003_sig000002c6
    );
  blk00000003_blk00000228 : XORCY
    port map (
      CI => blk00000003_sig000002d5,
      LI => blk00000003_sig000002d6,
      O => blk00000003_sig000002d7
    );
  blk00000003_blk00000227 : XORCY
    port map (
      CI => blk00000003_sig000002d2,
      LI => blk00000003_sig000002d3,
      O => blk00000003_sig000002d4
    );
  blk00000003_blk00000226 : XORCY
    port map (
      CI => blk00000003_sig000002cf,
      LI => blk00000003_sig000002d0,
      O => blk00000003_sig000002d1
    );
  blk00000003_blk00000225 : XORCY
    port map (
      CI => blk00000003_sig000002cc,
      LI => blk00000003_sig000002cd,
      O => blk00000003_sig000002ce
    );
  blk00000003_blk00000224 : XORCY
    port map (
      CI => blk00000003_sig000002c9,
      LI => blk00000003_sig000002ca,
      O => blk00000003_sig000002cb
    );
  blk00000003_blk00000223 : XORCY
    port map (
      CI => blk00000003_sig000002c6,
      LI => blk00000003_sig000002c7,
      O => blk00000003_sig000002c8
    );
  blk00000003_blk00000222 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002bc,
      Q => blk00000003_sig000002c5
    );
  blk00000003_blk00000221 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002ac,
      Q => blk00000003_sig000002c4
    );
  blk00000003_blk00000220 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002af,
      Q => blk00000003_sig000002c3
    );
  blk00000003_blk0000021f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002b2,
      Q => blk00000003_sig000002c2
    );
  blk00000003_blk0000021e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002b5,
      Q => blk00000003_sig000002c1
    );
  blk00000003_blk0000021d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002b8,
      Q => blk00000003_sig000002c0
    );
  blk00000003_blk0000021c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002bb,
      Q => blk00000003_sig000002bf
    );
  blk00000003_blk0000021b : MUXCY
    port map (
      CI => blk00000003_sig000002bd,
      DI => blk00000003_sig00000031,
      S => blk00000003_sig000002be,
      O => blk00000003_sig000002b9
    );
  blk00000003_blk0000021a : XORCY
    port map (
      CI => blk00000003_sig000002bd,
      LI => blk00000003_sig000002be,
      O => NLW_blk00000003_blk0000021a_O_UNCONNECTED
    );
  blk00000003_blk00000219 : MUXCY
    port map (
      CI => blk00000003_sig000002aa,
      DI => blk00000003_sig000002a7,
      S => blk00000003_sig000002ab,
      O => blk00000003_sig000002bc
    );
  blk00000003_blk00000218 : MUXCY
    port map (
      CI => blk00000003_sig000002b9,
      DI => blk00000003_sig000000c7,
      S => blk00000003_sig000002ba,
      O => blk00000003_sig000002b6
    );
  blk00000003_blk00000217 : MUXCY
    port map (
      CI => blk00000003_sig000002b6,
      DI => blk00000003_sig000002a3,
      S => blk00000003_sig000002b7,
      O => blk00000003_sig000002b3
    );
  blk00000003_blk00000216 : MUXCY
    port map (
      CI => blk00000003_sig000002b3,
      DI => blk00000003_sig000002a4,
      S => blk00000003_sig000002b4,
      O => blk00000003_sig000002b0
    );
  blk00000003_blk00000215 : MUXCY
    port map (
      CI => blk00000003_sig000002b0,
      DI => blk00000003_sig000002a5,
      S => blk00000003_sig000002b1,
      O => blk00000003_sig000002ad
    );
  blk00000003_blk00000214 : MUXCY
    port map (
      CI => blk00000003_sig000002ad,
      DI => blk00000003_sig000002a6,
      S => blk00000003_sig000002ae,
      O => blk00000003_sig000002aa
    );
  blk00000003_blk00000213 : XORCY
    port map (
      CI => blk00000003_sig000002b9,
      LI => blk00000003_sig000002ba,
      O => blk00000003_sig000002bb
    );
  blk00000003_blk00000212 : XORCY
    port map (
      CI => blk00000003_sig000002b6,
      LI => blk00000003_sig000002b7,
      O => blk00000003_sig000002b8
    );
  blk00000003_blk00000211 : XORCY
    port map (
      CI => blk00000003_sig000002b3,
      LI => blk00000003_sig000002b4,
      O => blk00000003_sig000002b5
    );
  blk00000003_blk00000210 : XORCY
    port map (
      CI => blk00000003_sig000002b0,
      LI => blk00000003_sig000002b1,
      O => blk00000003_sig000002b2
    );
  blk00000003_blk0000020f : XORCY
    port map (
      CI => blk00000003_sig000002ad,
      LI => blk00000003_sig000002ae,
      O => blk00000003_sig000002af
    );
  blk00000003_blk0000020e : XORCY
    port map (
      CI => blk00000003_sig000002aa,
      LI => blk00000003_sig000002ab,
      O => blk00000003_sig000002ac
    );
  blk00000003_blk0000020d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002a0,
      Q => blk00000003_sig000002a9
    );
  blk00000003_blk0000020c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000290,
      Q => blk00000003_sig000002a8
    );
  blk00000003_blk0000020b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000293,
      Q => blk00000003_sig000002a7
    );
  blk00000003_blk0000020a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000296,
      Q => blk00000003_sig000002a6
    );
  blk00000003_blk00000209 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000299,
      Q => blk00000003_sig000002a5
    );
  blk00000003_blk00000208 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000029c,
      Q => blk00000003_sig000002a4
    );
  blk00000003_blk00000207 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000029f,
      Q => blk00000003_sig000002a3
    );
  blk00000003_blk00000206 : MUXCY
    port map (
      CI => blk00000003_sig000002a1,
      DI => blk00000003_sig00000031,
      S => blk00000003_sig000002a2,
      O => blk00000003_sig0000029d
    );
  blk00000003_blk00000205 : XORCY
    port map (
      CI => blk00000003_sig000002a1,
      LI => blk00000003_sig000002a2,
      O => NLW_blk00000003_blk00000205_O_UNCONNECTED
    );
  blk00000003_blk00000204 : MUXCY
    port map (
      CI => blk00000003_sig0000028e,
      DI => blk00000003_sig0000028b,
      S => blk00000003_sig0000028f,
      O => blk00000003_sig000002a0
    );
  blk00000003_blk00000203 : MUXCY
    port map (
      CI => blk00000003_sig0000029d,
      DI => blk00000003_sig00000286,
      S => blk00000003_sig0000029e,
      O => blk00000003_sig0000029a
    );
  blk00000003_blk00000202 : MUXCY
    port map (
      CI => blk00000003_sig0000029a,
      DI => blk00000003_sig00000287,
      S => blk00000003_sig0000029b,
      O => blk00000003_sig00000297
    );
  blk00000003_blk00000201 : MUXCY
    port map (
      CI => blk00000003_sig00000297,
      DI => blk00000003_sig00000288,
      S => blk00000003_sig00000298,
      O => blk00000003_sig00000294
    );
  blk00000003_blk00000200 : MUXCY
    port map (
      CI => blk00000003_sig00000294,
      DI => blk00000003_sig00000289,
      S => blk00000003_sig00000295,
      O => blk00000003_sig00000291
    );
  blk00000003_blk000001ff : MUXCY
    port map (
      CI => blk00000003_sig00000291,
      DI => blk00000003_sig0000028a,
      S => blk00000003_sig00000292,
      O => blk00000003_sig0000028e
    );
  blk00000003_blk000001fe : XORCY
    port map (
      CI => blk00000003_sig0000029d,
      LI => blk00000003_sig0000029e,
      O => blk00000003_sig0000029f
    );
  blk00000003_blk000001fd : XORCY
    port map (
      CI => blk00000003_sig0000029a,
      LI => blk00000003_sig0000029b,
      O => blk00000003_sig0000029c
    );
  blk00000003_blk000001fc : XORCY
    port map (
      CI => blk00000003_sig00000297,
      LI => blk00000003_sig00000298,
      O => blk00000003_sig00000299
    );
  blk00000003_blk000001fb : XORCY
    port map (
      CI => blk00000003_sig00000294,
      LI => blk00000003_sig00000295,
      O => blk00000003_sig00000296
    );
  blk00000003_blk000001fa : XORCY
    port map (
      CI => blk00000003_sig00000291,
      LI => blk00000003_sig00000292,
      O => blk00000003_sig00000293
    );
  blk00000003_blk000001f9 : XORCY
    port map (
      CI => blk00000003_sig0000028e,
      LI => blk00000003_sig0000028f,
      O => blk00000003_sig00000290
    );
  blk00000003_blk000001f8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000282,
      Q => blk00000003_sig0000028d
    );
  blk00000003_blk000001f7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000272,
      Q => blk00000003_sig0000028c
    );
  blk00000003_blk000001f6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000275,
      Q => blk00000003_sig0000028b
    );
  blk00000003_blk000001f5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000278,
      Q => blk00000003_sig0000028a
    );
  blk00000003_blk000001f4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000027b,
      Q => blk00000003_sig00000289
    );
  blk00000003_blk000001f3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000027e,
      Q => blk00000003_sig00000288
    );
  blk00000003_blk000001f2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000281,
      Q => blk00000003_sig00000287
    );
  blk00000003_blk000001f1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000285,
      Q => blk00000003_sig00000286
    );
  blk00000003_blk000001f0 : MUXCY
    port map (
      CI => blk00000003_sig00000283,
      DI => blk00000003_sig00000078,
      S => blk00000003_sig00000284,
      O => blk00000003_sig0000027f
    );
  blk00000003_blk000001ef : XORCY
    port map (
      CI => blk00000003_sig00000283,
      LI => blk00000003_sig00000284,
      O => blk00000003_sig00000285
    );
  blk00000003_blk000001ee : MUXCY
    port map (
      CI => blk00000003_sig00000270,
      DI => blk00000003_sig0000026d,
      S => blk00000003_sig00000271,
      O => blk00000003_sig00000282
    );
  blk00000003_blk000001ed : MUXCY
    port map (
      CI => blk00000003_sig0000027f,
      DI => blk00000003_sig00000268,
      S => blk00000003_sig00000280,
      O => blk00000003_sig0000027c
    );
  blk00000003_blk000001ec : MUXCY
    port map (
      CI => blk00000003_sig0000027c,
      DI => blk00000003_sig00000269,
      S => blk00000003_sig0000027d,
      O => blk00000003_sig00000279
    );
  blk00000003_blk000001eb : MUXCY
    port map (
      CI => blk00000003_sig00000279,
      DI => blk00000003_sig0000026a,
      S => blk00000003_sig0000027a,
      O => blk00000003_sig00000276
    );
  blk00000003_blk000001ea : MUXCY
    port map (
      CI => blk00000003_sig00000276,
      DI => blk00000003_sig0000026b,
      S => blk00000003_sig00000277,
      O => blk00000003_sig00000273
    );
  blk00000003_blk000001e9 : MUXCY
    port map (
      CI => blk00000003_sig00000273,
      DI => blk00000003_sig0000026c,
      S => blk00000003_sig00000274,
      O => blk00000003_sig00000270
    );
  blk00000003_blk000001e8 : XORCY
    port map (
      CI => blk00000003_sig0000027f,
      LI => blk00000003_sig00000280,
      O => blk00000003_sig00000281
    );
  blk00000003_blk000001e7 : XORCY
    port map (
      CI => blk00000003_sig0000027c,
      LI => blk00000003_sig0000027d,
      O => blk00000003_sig0000027e
    );
  blk00000003_blk000001e6 : XORCY
    port map (
      CI => blk00000003_sig00000279,
      LI => blk00000003_sig0000027a,
      O => blk00000003_sig0000027b
    );
  blk00000003_blk000001e5 : XORCY
    port map (
      CI => blk00000003_sig00000276,
      LI => blk00000003_sig00000277,
      O => blk00000003_sig00000278
    );
  blk00000003_blk000001e4 : XORCY
    port map (
      CI => blk00000003_sig00000273,
      LI => blk00000003_sig00000274,
      O => blk00000003_sig00000275
    );
  blk00000003_blk000001e3 : XORCY
    port map (
      CI => blk00000003_sig00000270,
      LI => blk00000003_sig00000271,
      O => blk00000003_sig00000272
    );
  blk00000003_blk000001e2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000264,
      Q => blk00000003_sig0000026f
    );
  blk00000003_blk000001e1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000254,
      Q => blk00000003_sig0000026e
    );
  blk00000003_blk000001e0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000257,
      Q => blk00000003_sig0000026d
    );
  blk00000003_blk000001df : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000025a,
      Q => blk00000003_sig0000026c
    );
  blk00000003_blk000001de : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000025d,
      Q => blk00000003_sig0000026b
    );
  blk00000003_blk000001dd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000260,
      Q => blk00000003_sig0000026a
    );
  blk00000003_blk000001dc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000263,
      Q => blk00000003_sig00000269
    );
  blk00000003_blk000001db : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000267,
      Q => blk00000003_sig00000268
    );
  blk00000003_blk000001da : MUXCY
    port map (
      CI => blk00000003_sig00000265,
      DI => blk00000003_sig00000036,
      S => blk00000003_sig00000266,
      O => blk00000003_sig00000261
    );
  blk00000003_blk000001d9 : XORCY
    port map (
      CI => blk00000003_sig00000265,
      LI => blk00000003_sig00000266,
      O => blk00000003_sig00000267
    );
  blk00000003_blk000001d8 : MUXCY
    port map (
      CI => blk00000003_sig00000252,
      DI => blk00000003_sig0000024f,
      S => blk00000003_sig00000253,
      O => blk00000003_sig00000264
    );
  blk00000003_blk000001d7 : MUXCY
    port map (
      CI => blk00000003_sig00000261,
      DI => blk00000003_sig0000024a,
      S => blk00000003_sig00000262,
      O => blk00000003_sig0000025e
    );
  blk00000003_blk000001d6 : MUXCY
    port map (
      CI => blk00000003_sig0000025e,
      DI => blk00000003_sig0000024b,
      S => blk00000003_sig0000025f,
      O => blk00000003_sig0000025b
    );
  blk00000003_blk000001d5 : MUXCY
    port map (
      CI => blk00000003_sig0000025b,
      DI => blk00000003_sig0000024c,
      S => blk00000003_sig0000025c,
      O => blk00000003_sig00000258
    );
  blk00000003_blk000001d4 : MUXCY
    port map (
      CI => blk00000003_sig00000258,
      DI => blk00000003_sig0000024d,
      S => blk00000003_sig00000259,
      O => blk00000003_sig00000255
    );
  blk00000003_blk000001d3 : MUXCY
    port map (
      CI => blk00000003_sig00000255,
      DI => blk00000003_sig0000024e,
      S => blk00000003_sig00000256,
      O => blk00000003_sig00000252
    );
  blk00000003_blk000001d2 : XORCY
    port map (
      CI => blk00000003_sig00000261,
      LI => blk00000003_sig00000262,
      O => blk00000003_sig00000263
    );
  blk00000003_blk000001d1 : XORCY
    port map (
      CI => blk00000003_sig0000025e,
      LI => blk00000003_sig0000025f,
      O => blk00000003_sig00000260
    );
  blk00000003_blk000001d0 : XORCY
    port map (
      CI => blk00000003_sig0000025b,
      LI => blk00000003_sig0000025c,
      O => blk00000003_sig0000025d
    );
  blk00000003_blk000001cf : XORCY
    port map (
      CI => blk00000003_sig00000258,
      LI => blk00000003_sig00000259,
      O => blk00000003_sig0000025a
    );
  blk00000003_blk000001ce : XORCY
    port map (
      CI => blk00000003_sig00000255,
      LI => blk00000003_sig00000256,
      O => blk00000003_sig00000257
    );
  blk00000003_blk000001cd : XORCY
    port map (
      CI => blk00000003_sig00000252,
      LI => blk00000003_sig00000253,
      O => blk00000003_sig00000254
    );
  blk00000003_blk000001cc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000246,
      Q => blk00000003_sig00000251
    );
  blk00000003_blk000001cb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000236,
      Q => blk00000003_sig00000250
    );
  blk00000003_blk000001ca : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000239,
      Q => blk00000003_sig0000024f
    );
  blk00000003_blk000001c9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000023c,
      Q => blk00000003_sig0000024e
    );
  blk00000003_blk000001c8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000023f,
      Q => blk00000003_sig0000024d
    );
  blk00000003_blk000001c7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000242,
      Q => blk00000003_sig0000024c
    );
  blk00000003_blk000001c6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000245,
      Q => blk00000003_sig0000024b
    );
  blk00000003_blk000001c5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000249,
      Q => blk00000003_sig0000024a
    );
  blk00000003_blk000001c4 : MUXCY
    port map (
      CI => blk00000003_sig00000247,
      DI => blk00000003_sig0000003a,
      S => blk00000003_sig00000248,
      O => blk00000003_sig00000243
    );
  blk00000003_blk000001c3 : XORCY
    port map (
      CI => blk00000003_sig00000247,
      LI => blk00000003_sig00000248,
      O => blk00000003_sig00000249
    );
  blk00000003_blk000001c2 : MUXCY
    port map (
      CI => blk00000003_sig00000234,
      DI => blk00000003_sig00000231,
      S => blk00000003_sig00000235,
      O => blk00000003_sig00000246
    );
  blk00000003_blk000001c1 : MUXCY
    port map (
      CI => blk00000003_sig00000243,
      DI => blk00000003_sig0000022c,
      S => blk00000003_sig00000244,
      O => blk00000003_sig00000240
    );
  blk00000003_blk000001c0 : MUXCY
    port map (
      CI => blk00000003_sig00000240,
      DI => blk00000003_sig0000022d,
      S => blk00000003_sig00000241,
      O => blk00000003_sig0000023d
    );
  blk00000003_blk000001bf : MUXCY
    port map (
      CI => blk00000003_sig0000023d,
      DI => blk00000003_sig0000022e,
      S => blk00000003_sig0000023e,
      O => blk00000003_sig0000023a
    );
  blk00000003_blk000001be : MUXCY
    port map (
      CI => blk00000003_sig0000023a,
      DI => blk00000003_sig0000022f,
      S => blk00000003_sig0000023b,
      O => blk00000003_sig00000237
    );
  blk00000003_blk000001bd : MUXCY
    port map (
      CI => blk00000003_sig00000237,
      DI => blk00000003_sig00000230,
      S => blk00000003_sig00000238,
      O => blk00000003_sig00000234
    );
  blk00000003_blk000001bc : XORCY
    port map (
      CI => blk00000003_sig00000243,
      LI => blk00000003_sig00000244,
      O => blk00000003_sig00000245
    );
  blk00000003_blk000001bb : XORCY
    port map (
      CI => blk00000003_sig00000240,
      LI => blk00000003_sig00000241,
      O => blk00000003_sig00000242
    );
  blk00000003_blk000001ba : XORCY
    port map (
      CI => blk00000003_sig0000023d,
      LI => blk00000003_sig0000023e,
      O => blk00000003_sig0000023f
    );
  blk00000003_blk000001b9 : XORCY
    port map (
      CI => blk00000003_sig0000023a,
      LI => blk00000003_sig0000023b,
      O => blk00000003_sig0000023c
    );
  blk00000003_blk000001b8 : XORCY
    port map (
      CI => blk00000003_sig00000237,
      LI => blk00000003_sig00000238,
      O => blk00000003_sig00000239
    );
  blk00000003_blk000001b7 : XORCY
    port map (
      CI => blk00000003_sig00000234,
      LI => blk00000003_sig00000235,
      O => blk00000003_sig00000236
    );
  blk00000003_blk000001b6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000228,
      Q => blk00000003_sig00000233
    );
  blk00000003_blk000001b5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000218,
      Q => blk00000003_sig00000232
    );
  blk00000003_blk000001b4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000021b,
      Q => blk00000003_sig00000231
    );
  blk00000003_blk000001b3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000021e,
      Q => blk00000003_sig00000230
    );
  blk00000003_blk000001b2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000221,
      Q => blk00000003_sig0000022f
    );
  blk00000003_blk000001b1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000224,
      Q => blk00000003_sig0000022e
    );
  blk00000003_blk000001b0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000227,
      Q => blk00000003_sig0000022d
    );
  blk00000003_blk000001af : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000022b,
      Q => blk00000003_sig0000022c
    );
  blk00000003_blk000001ae : MUXCY
    port map (
      CI => blk00000003_sig00000229,
      DI => blk00000003_sig0000003f,
      S => blk00000003_sig0000022a,
      O => blk00000003_sig00000225
    );
  blk00000003_blk000001ad : XORCY
    port map (
      CI => blk00000003_sig00000229,
      LI => blk00000003_sig0000022a,
      O => blk00000003_sig0000022b
    );
  blk00000003_blk000001ac : MUXCY
    port map (
      CI => blk00000003_sig00000216,
      DI => blk00000003_sig00000213,
      S => blk00000003_sig00000217,
      O => blk00000003_sig00000228
    );
  blk00000003_blk000001ab : MUXCY
    port map (
      CI => blk00000003_sig00000225,
      DI => blk00000003_sig0000020e,
      S => blk00000003_sig00000226,
      O => blk00000003_sig00000222
    );
  blk00000003_blk000001aa : MUXCY
    port map (
      CI => blk00000003_sig00000222,
      DI => blk00000003_sig0000020f,
      S => blk00000003_sig00000223,
      O => blk00000003_sig0000021f
    );
  blk00000003_blk000001a9 : MUXCY
    port map (
      CI => blk00000003_sig0000021f,
      DI => blk00000003_sig00000210,
      S => blk00000003_sig00000220,
      O => blk00000003_sig0000021c
    );
  blk00000003_blk000001a8 : MUXCY
    port map (
      CI => blk00000003_sig0000021c,
      DI => blk00000003_sig00000211,
      S => blk00000003_sig0000021d,
      O => blk00000003_sig00000219
    );
  blk00000003_blk000001a7 : MUXCY
    port map (
      CI => blk00000003_sig00000219,
      DI => blk00000003_sig00000212,
      S => blk00000003_sig0000021a,
      O => blk00000003_sig00000216
    );
  blk00000003_blk000001a6 : XORCY
    port map (
      CI => blk00000003_sig00000225,
      LI => blk00000003_sig00000226,
      O => blk00000003_sig00000227
    );
  blk00000003_blk000001a5 : XORCY
    port map (
      CI => blk00000003_sig00000222,
      LI => blk00000003_sig00000223,
      O => blk00000003_sig00000224
    );
  blk00000003_blk000001a4 : XORCY
    port map (
      CI => blk00000003_sig0000021f,
      LI => blk00000003_sig00000220,
      O => blk00000003_sig00000221
    );
  blk00000003_blk000001a3 : XORCY
    port map (
      CI => blk00000003_sig0000021c,
      LI => blk00000003_sig0000021d,
      O => blk00000003_sig0000021e
    );
  blk00000003_blk000001a2 : XORCY
    port map (
      CI => blk00000003_sig00000219,
      LI => blk00000003_sig0000021a,
      O => blk00000003_sig0000021b
    );
  blk00000003_blk000001a1 : XORCY
    port map (
      CI => blk00000003_sig00000216,
      LI => blk00000003_sig00000217,
      O => blk00000003_sig00000218
    );
  blk00000003_blk000001a0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000020a,
      Q => blk00000003_sig00000215
    );
  blk00000003_blk0000019f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001fa,
      Q => blk00000003_sig00000214
    );
  blk00000003_blk0000019e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001fd,
      Q => blk00000003_sig00000213
    );
  blk00000003_blk0000019d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000200,
      Q => blk00000003_sig00000212
    );
  blk00000003_blk0000019c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000203,
      Q => blk00000003_sig00000211
    );
  blk00000003_blk0000019b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000206,
      Q => blk00000003_sig00000210
    );
  blk00000003_blk0000019a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000209,
      Q => blk00000003_sig0000020f
    );
  blk00000003_blk00000199 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000020d,
      Q => blk00000003_sig0000020e
    );
  blk00000003_blk00000198 : MUXCY
    port map (
      CI => blk00000003_sig0000020b,
      DI => blk00000003_sig00000045,
      S => blk00000003_sig0000020c,
      O => blk00000003_sig00000207
    );
  blk00000003_blk00000197 : XORCY
    port map (
      CI => blk00000003_sig0000020b,
      LI => blk00000003_sig0000020c,
      O => blk00000003_sig0000020d
    );
  blk00000003_blk00000196 : MUXCY
    port map (
      CI => blk00000003_sig000001f8,
      DI => blk00000003_sig000001f6,
      S => blk00000003_sig000001f9,
      O => blk00000003_sig0000020a
    );
  blk00000003_blk00000195 : MUXCY
    port map (
      CI => blk00000003_sig00000207,
      DI => blk00000003_sig000001f1,
      S => blk00000003_sig00000208,
      O => blk00000003_sig00000204
    );
  blk00000003_blk00000194 : MUXCY
    port map (
      CI => blk00000003_sig00000204,
      DI => blk00000003_sig000001f2,
      S => blk00000003_sig00000205,
      O => blk00000003_sig00000201
    );
  blk00000003_blk00000193 : MUXCY
    port map (
      CI => blk00000003_sig00000201,
      DI => blk00000003_sig000001f3,
      S => blk00000003_sig00000202,
      O => blk00000003_sig000001fe
    );
  blk00000003_blk00000192 : MUXCY
    port map (
      CI => blk00000003_sig000001fe,
      DI => blk00000003_sig000001f4,
      S => blk00000003_sig000001ff,
      O => blk00000003_sig000001fb
    );
  blk00000003_blk00000191 : MUXCY
    port map (
      CI => blk00000003_sig000001fb,
      DI => blk00000003_sig000001f5,
      S => blk00000003_sig000001fc,
      O => blk00000003_sig000001f8
    );
  blk00000003_blk00000190 : XORCY
    port map (
      CI => blk00000003_sig00000207,
      LI => blk00000003_sig00000208,
      O => blk00000003_sig00000209
    );
  blk00000003_blk0000018f : XORCY
    port map (
      CI => blk00000003_sig00000204,
      LI => blk00000003_sig00000205,
      O => blk00000003_sig00000206
    );
  blk00000003_blk0000018e : XORCY
    port map (
      CI => blk00000003_sig00000201,
      LI => blk00000003_sig00000202,
      O => blk00000003_sig00000203
    );
  blk00000003_blk0000018d : XORCY
    port map (
      CI => blk00000003_sig000001fe,
      LI => blk00000003_sig000001ff,
      O => blk00000003_sig00000200
    );
  blk00000003_blk0000018c : XORCY
    port map (
      CI => blk00000003_sig000001fb,
      LI => blk00000003_sig000001fc,
      O => blk00000003_sig000001fd
    );
  blk00000003_blk0000018b : XORCY
    port map (
      CI => blk00000003_sig000001f8,
      LI => blk00000003_sig000001f9,
      O => blk00000003_sig000001fa
    );
  blk00000003_blk0000018a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001ed,
      Q => blk00000003_sig000001f7
    );
  blk00000003_blk00000189 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001dd,
      Q => blk00000003_sig00000070
    );
  blk00000003_blk00000188 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001e0,
      Q => blk00000003_sig000001f6
    );
  blk00000003_blk00000187 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001e3,
      Q => blk00000003_sig000001f5
    );
  blk00000003_blk00000186 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001e6,
      Q => blk00000003_sig000001f4
    );
  blk00000003_blk00000185 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001e9,
      Q => blk00000003_sig000001f3
    );
  blk00000003_blk00000184 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001ec,
      Q => blk00000003_sig000001f2
    );
  blk00000003_blk00000183 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001f0,
      Q => blk00000003_sig000001f1
    );
  blk00000003_blk00000182 : MUXCY
    port map (
      CI => blk00000003_sig000001ee,
      DI => blk00000003_sig00000058,
      S => blk00000003_sig000001ef,
      O => blk00000003_sig000001ea
    );
  blk00000003_blk00000181 : XORCY
    port map (
      CI => blk00000003_sig000001ee,
      LI => blk00000003_sig000001ef,
      O => blk00000003_sig000001f0
    );
  blk00000003_blk00000180 : MUXCY
    port map (
      CI => blk00000003_sig000001db,
      DI => blk00000003_sig000001d9,
      S => blk00000003_sig000001dc,
      O => blk00000003_sig000001ed
    );
  blk00000003_blk0000017f : MUXCY
    port map (
      CI => blk00000003_sig000001ea,
      DI => blk00000003_sig000001d4,
      S => blk00000003_sig000001eb,
      O => blk00000003_sig000001e7
    );
  blk00000003_blk0000017e : MUXCY
    port map (
      CI => blk00000003_sig000001e7,
      DI => blk00000003_sig000001d5,
      S => blk00000003_sig000001e8,
      O => blk00000003_sig000001e4
    );
  blk00000003_blk0000017d : MUXCY
    port map (
      CI => blk00000003_sig000001e4,
      DI => blk00000003_sig000001d6,
      S => blk00000003_sig000001e5,
      O => blk00000003_sig000001e1
    );
  blk00000003_blk0000017c : MUXCY
    port map (
      CI => blk00000003_sig000001e1,
      DI => blk00000003_sig000001d7,
      S => blk00000003_sig000001e2,
      O => blk00000003_sig000001de
    );
  blk00000003_blk0000017b : MUXCY
    port map (
      CI => blk00000003_sig000001de,
      DI => blk00000003_sig000001d8,
      S => blk00000003_sig000001df,
      O => blk00000003_sig000001db
    );
  blk00000003_blk0000017a : XORCY
    port map (
      CI => blk00000003_sig000001ea,
      LI => blk00000003_sig000001eb,
      O => blk00000003_sig000001ec
    );
  blk00000003_blk00000179 : XORCY
    port map (
      CI => blk00000003_sig000001e7,
      LI => blk00000003_sig000001e8,
      O => blk00000003_sig000001e9
    );
  blk00000003_blk00000178 : XORCY
    port map (
      CI => blk00000003_sig000001e4,
      LI => blk00000003_sig000001e5,
      O => blk00000003_sig000001e6
    );
  blk00000003_blk00000177 : XORCY
    port map (
      CI => blk00000003_sig000001e1,
      LI => blk00000003_sig000001e2,
      O => blk00000003_sig000001e3
    );
  blk00000003_blk00000176 : XORCY
    port map (
      CI => blk00000003_sig000001de,
      LI => blk00000003_sig000001df,
      O => blk00000003_sig000001e0
    );
  blk00000003_blk00000175 : XORCY
    port map (
      CI => blk00000003_sig000001db,
      LI => blk00000003_sig000001dc,
      O => blk00000003_sig000001dd
    );
  blk00000003_blk00000174 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001d0,
      Q => blk00000003_sig000001da
    );
  blk00000003_blk00000173 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001c0,
      Q => blk00000003_sig00000046
    );
  blk00000003_blk00000172 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001c3,
      Q => blk00000003_sig000001d9
    );
  blk00000003_blk00000171 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001c6,
      Q => blk00000003_sig000001d8
    );
  blk00000003_blk00000170 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001c9,
      Q => blk00000003_sig000001d7
    );
  blk00000003_blk0000016f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001cc,
      Q => blk00000003_sig000001d6
    );
  blk00000003_blk0000016e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001cf,
      Q => blk00000003_sig000001d5
    );
  blk00000003_blk0000016d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001d3,
      Q => blk00000003_sig000001d4
    );
  blk00000003_blk0000016c : MUXCY
    port map (
      CI => blk00000003_sig000001d1,
      DI => blk00000003_sig00000065,
      S => blk00000003_sig000001d2,
      O => blk00000003_sig000001cd
    );
  blk00000003_blk0000016b : XORCY
    port map (
      CI => blk00000003_sig000001d1,
      LI => blk00000003_sig000001d2,
      O => blk00000003_sig000001d3
    );
  blk00000003_blk0000016a : MUXCY
    port map (
      CI => blk00000003_sig000001be,
      DI => blk00000003_sig000001bc,
      S => blk00000003_sig000001bf,
      O => blk00000003_sig000001d0
    );
  blk00000003_blk00000169 : MUXCY
    port map (
      CI => blk00000003_sig000001cd,
      DI => blk00000003_sig000001b7,
      S => blk00000003_sig000001ce,
      O => blk00000003_sig000001ca
    );
  blk00000003_blk00000168 : MUXCY
    port map (
      CI => blk00000003_sig000001ca,
      DI => blk00000003_sig000001b8,
      S => blk00000003_sig000001cb,
      O => blk00000003_sig000001c7
    );
  blk00000003_blk00000167 : MUXCY
    port map (
      CI => blk00000003_sig000001c7,
      DI => blk00000003_sig000001b9,
      S => blk00000003_sig000001c8,
      O => blk00000003_sig000001c4
    );
  blk00000003_blk00000166 : MUXCY
    port map (
      CI => blk00000003_sig000001c4,
      DI => blk00000003_sig000001ba,
      S => blk00000003_sig000001c5,
      O => blk00000003_sig000001c1
    );
  blk00000003_blk00000165 : MUXCY
    port map (
      CI => blk00000003_sig000001c1,
      DI => blk00000003_sig000001bb,
      S => blk00000003_sig000001c2,
      O => blk00000003_sig000001be
    );
  blk00000003_blk00000164 : XORCY
    port map (
      CI => blk00000003_sig000001cd,
      LI => blk00000003_sig000001ce,
      O => blk00000003_sig000001cf
    );
  blk00000003_blk00000163 : XORCY
    port map (
      CI => blk00000003_sig000001ca,
      LI => blk00000003_sig000001cb,
      O => blk00000003_sig000001cc
    );
  blk00000003_blk00000162 : XORCY
    port map (
      CI => blk00000003_sig000001c7,
      LI => blk00000003_sig000001c8,
      O => blk00000003_sig000001c9
    );
  blk00000003_blk00000161 : XORCY
    port map (
      CI => blk00000003_sig000001c4,
      LI => blk00000003_sig000001c5,
      O => blk00000003_sig000001c6
    );
  blk00000003_blk00000160 : XORCY
    port map (
      CI => blk00000003_sig000001c1,
      LI => blk00000003_sig000001c2,
      O => blk00000003_sig000001c3
    );
  blk00000003_blk0000015f : XORCY
    port map (
      CI => blk00000003_sig000001be,
      LI => blk00000003_sig000001bf,
      O => blk00000003_sig000001c0
    );
  blk00000003_blk0000015e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001b2,
      Q => blk00000003_sig000001bd
    );
  blk00000003_blk0000015d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001a2,
      Q => blk00000003_sig00000059
    );
  blk00000003_blk0000015c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001a5,
      Q => blk00000003_sig000001bc
    );
  blk00000003_blk0000015b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001a8,
      Q => blk00000003_sig000001bb
    );
  blk00000003_blk0000015a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001ab,
      Q => blk00000003_sig000001ba
    );
  blk00000003_blk00000159 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001ae,
      Q => blk00000003_sig000001b9
    );
  blk00000003_blk00000158 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001b1,
      Q => blk00000003_sig000001b8
    );
  blk00000003_blk00000157 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001b5,
      Q => blk00000003_sig000001b7
    );
  blk00000003_blk00000156 : MUXCY
    port map (
      CI => blk00000003_sig000001b3,
      DI => blk00000003_sig000001b6,
      S => blk00000003_sig000001b4,
      O => blk00000003_sig000001af
    );
  blk00000003_blk00000155 : XORCY
    port map (
      CI => blk00000003_sig000001b3,
      LI => blk00000003_sig000001b4,
      O => blk00000003_sig000001b5
    );
  blk00000003_blk00000154 : MUXCY
    port map (
      CI => blk00000003_sig000001a0,
      DI => blk00000003_sig0000019e,
      S => blk00000003_sig000001a1,
      O => blk00000003_sig000001b2
    );
  blk00000003_blk00000153 : MUXCY
    port map (
      CI => blk00000003_sig000001af,
      DI => blk00000003_sig00000199,
      S => blk00000003_sig000001b0,
      O => blk00000003_sig000001ac
    );
  blk00000003_blk00000152 : MUXCY
    port map (
      CI => blk00000003_sig000001ac,
      DI => blk00000003_sig0000019a,
      S => blk00000003_sig000001ad,
      O => blk00000003_sig000001a9
    );
  blk00000003_blk00000151 : MUXCY
    port map (
      CI => blk00000003_sig000001a9,
      DI => blk00000003_sig0000019b,
      S => blk00000003_sig000001aa,
      O => blk00000003_sig000001a6
    );
  blk00000003_blk00000150 : MUXCY
    port map (
      CI => blk00000003_sig000001a6,
      DI => blk00000003_sig0000019c,
      S => blk00000003_sig000001a7,
      O => blk00000003_sig000001a3
    );
  blk00000003_blk0000014f : MUXCY
    port map (
      CI => blk00000003_sig000001a3,
      DI => blk00000003_sig0000019d,
      S => blk00000003_sig000001a4,
      O => blk00000003_sig000001a0
    );
  blk00000003_blk0000014e : XORCY
    port map (
      CI => blk00000003_sig000001af,
      LI => blk00000003_sig000001b0,
      O => blk00000003_sig000001b1
    );
  blk00000003_blk0000014d : XORCY
    port map (
      CI => blk00000003_sig000001ac,
      LI => blk00000003_sig000001ad,
      O => blk00000003_sig000001ae
    );
  blk00000003_blk0000014c : XORCY
    port map (
      CI => blk00000003_sig000001a9,
      LI => blk00000003_sig000001aa,
      O => blk00000003_sig000001ab
    );
  blk00000003_blk0000014b : XORCY
    port map (
      CI => blk00000003_sig000001a6,
      LI => blk00000003_sig000001a7,
      O => blk00000003_sig000001a8
    );
  blk00000003_blk0000014a : XORCY
    port map (
      CI => blk00000003_sig000001a3,
      LI => blk00000003_sig000001a4,
      O => blk00000003_sig000001a5
    );
  blk00000003_blk00000149 : XORCY
    port map (
      CI => blk00000003_sig000001a0,
      LI => blk00000003_sig000001a1,
      O => blk00000003_sig000001a2
    );
  blk00000003_blk00000148 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000194,
      Q => blk00000003_sig0000019f
    );
  blk00000003_blk00000147 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000184,
      Q => blk00000003_sig00000066
    );
  blk00000003_blk00000146 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000187,
      Q => blk00000003_sig0000019e
    );
  blk00000003_blk00000145 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000018a,
      Q => blk00000003_sig0000019d
    );
  blk00000003_blk00000144 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000018d,
      Q => blk00000003_sig0000019c
    );
  blk00000003_blk00000143 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000190,
      Q => blk00000003_sig0000019b
    );
  blk00000003_blk00000142 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000193,
      Q => blk00000003_sig0000019a
    );
  blk00000003_blk00000141 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000197,
      Q => blk00000003_sig00000199
    );
  blk00000003_blk00000140 : MUXCY
    port map (
      CI => blk00000003_sig00000195,
      DI => blk00000003_sig00000198,
      S => blk00000003_sig00000196,
      O => blk00000003_sig00000191
    );
  blk00000003_blk0000013f : XORCY
    port map (
      CI => blk00000003_sig00000195,
      LI => blk00000003_sig00000196,
      O => blk00000003_sig00000197
    );
  blk00000003_blk0000013e : MUXCY
    port map (
      CI => blk00000003_sig00000182,
      DI => blk00000003_sig00000180,
      S => blk00000003_sig00000183,
      O => blk00000003_sig00000194
    );
  blk00000003_blk0000013d : MUXCY
    port map (
      CI => blk00000003_sig00000191,
      DI => blk00000003_sig0000017b,
      S => blk00000003_sig00000192,
      O => blk00000003_sig0000018e
    );
  blk00000003_blk0000013c : MUXCY
    port map (
      CI => blk00000003_sig0000018e,
      DI => blk00000003_sig0000017c,
      S => blk00000003_sig0000018f,
      O => blk00000003_sig0000018b
    );
  blk00000003_blk0000013b : MUXCY
    port map (
      CI => blk00000003_sig0000018b,
      DI => blk00000003_sig0000017d,
      S => blk00000003_sig0000018c,
      O => blk00000003_sig00000188
    );
  blk00000003_blk0000013a : MUXCY
    port map (
      CI => blk00000003_sig00000188,
      DI => blk00000003_sig0000017e,
      S => blk00000003_sig00000189,
      O => blk00000003_sig00000185
    );
  blk00000003_blk00000139 : MUXCY
    port map (
      CI => blk00000003_sig00000185,
      DI => blk00000003_sig0000017f,
      S => blk00000003_sig00000186,
      O => blk00000003_sig00000182
    );
  blk00000003_blk00000138 : XORCY
    port map (
      CI => blk00000003_sig00000191,
      LI => blk00000003_sig00000192,
      O => blk00000003_sig00000193
    );
  blk00000003_blk00000137 : XORCY
    port map (
      CI => blk00000003_sig0000018e,
      LI => blk00000003_sig0000018f,
      O => blk00000003_sig00000190
    );
  blk00000003_blk00000136 : XORCY
    port map (
      CI => blk00000003_sig0000018b,
      LI => blk00000003_sig0000018c,
      O => blk00000003_sig0000018d
    );
  blk00000003_blk00000135 : XORCY
    port map (
      CI => blk00000003_sig00000188,
      LI => blk00000003_sig00000189,
      O => blk00000003_sig0000018a
    );
  blk00000003_blk00000134 : XORCY
    port map (
      CI => blk00000003_sig00000185,
      LI => blk00000003_sig00000186,
      O => blk00000003_sig00000187
    );
  blk00000003_blk00000133 : XORCY
    port map (
      CI => blk00000003_sig00000182,
      LI => blk00000003_sig00000183,
      O => blk00000003_sig00000184
    );
  blk00000003_blk00000132 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000176,
      Q => blk00000003_sig00000181
    );
  blk00000003_blk00000131 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000166,
      Q => blk00000003_sig0000006a
    );
  blk00000003_blk00000130 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000169,
      Q => blk00000003_sig00000180
    );
  blk00000003_blk0000012f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000016c,
      Q => blk00000003_sig0000017f
    );
  blk00000003_blk0000012e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000016f,
      Q => blk00000003_sig0000017e
    );
  blk00000003_blk0000012d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000172,
      Q => blk00000003_sig0000017d
    );
  blk00000003_blk0000012c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000175,
      Q => blk00000003_sig0000017c
    );
  blk00000003_blk0000012b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000179,
      Q => blk00000003_sig0000017b
    );
  blk00000003_blk0000012a : MUXCY
    port map (
      CI => blk00000003_sig00000177,
      DI => blk00000003_sig0000017a,
      S => blk00000003_sig00000178,
      O => blk00000003_sig00000173
    );
  blk00000003_blk00000129 : XORCY
    port map (
      CI => blk00000003_sig00000177,
      LI => blk00000003_sig00000178,
      O => blk00000003_sig00000179
    );
  blk00000003_blk00000128 : MUXCY
    port map (
      CI => blk00000003_sig00000164,
      DI => blk00000003_sig00000162,
      S => blk00000003_sig00000165,
      O => blk00000003_sig00000176
    );
  blk00000003_blk00000127 : MUXCY
    port map (
      CI => blk00000003_sig00000173,
      DI => blk00000003_sig0000015d,
      S => blk00000003_sig00000174,
      O => blk00000003_sig00000170
    );
  blk00000003_blk00000126 : MUXCY
    port map (
      CI => blk00000003_sig00000170,
      DI => blk00000003_sig0000015e,
      S => blk00000003_sig00000171,
      O => blk00000003_sig0000016d
    );
  blk00000003_blk00000125 : MUXCY
    port map (
      CI => blk00000003_sig0000016d,
      DI => blk00000003_sig0000015f,
      S => blk00000003_sig0000016e,
      O => blk00000003_sig0000016a
    );
  blk00000003_blk00000124 : MUXCY
    port map (
      CI => blk00000003_sig0000016a,
      DI => blk00000003_sig00000160,
      S => blk00000003_sig0000016b,
      O => blk00000003_sig00000167
    );
  blk00000003_blk00000123 : MUXCY
    port map (
      CI => blk00000003_sig00000167,
      DI => blk00000003_sig00000161,
      S => blk00000003_sig00000168,
      O => blk00000003_sig00000164
    );
  blk00000003_blk00000122 : XORCY
    port map (
      CI => blk00000003_sig00000173,
      LI => blk00000003_sig00000174,
      O => blk00000003_sig00000175
    );
  blk00000003_blk00000121 : XORCY
    port map (
      CI => blk00000003_sig00000170,
      LI => blk00000003_sig00000171,
      O => blk00000003_sig00000172
    );
  blk00000003_blk00000120 : XORCY
    port map (
      CI => blk00000003_sig0000016d,
      LI => blk00000003_sig0000016e,
      O => blk00000003_sig0000016f
    );
  blk00000003_blk0000011f : XORCY
    port map (
      CI => blk00000003_sig0000016a,
      LI => blk00000003_sig0000016b,
      O => blk00000003_sig0000016c
    );
  blk00000003_blk0000011e : XORCY
    port map (
      CI => blk00000003_sig00000167,
      LI => blk00000003_sig00000168,
      O => blk00000003_sig00000169
    );
  blk00000003_blk0000011d : XORCY
    port map (
      CI => blk00000003_sig00000164,
      LI => blk00000003_sig00000165,
      O => blk00000003_sig00000166
    );
  blk00000003_blk0000011c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000158,
      Q => blk00000003_sig00000163
    );
  blk00000003_blk0000011b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000148,
      Q => blk00000003_sig0000006d
    );
  blk00000003_blk0000011a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000014b,
      Q => blk00000003_sig00000162
    );
  blk00000003_blk00000119 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000014e,
      Q => blk00000003_sig00000161
    );
  blk00000003_blk00000118 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000151,
      Q => blk00000003_sig00000160
    );
  blk00000003_blk00000117 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000154,
      Q => blk00000003_sig0000015f
    );
  blk00000003_blk00000116 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000157,
      Q => blk00000003_sig0000015e
    );
  blk00000003_blk00000115 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000015b,
      Q => blk00000003_sig0000015d
    );
  blk00000003_blk00000114 : MUXCY
    port map (
      CI => blk00000003_sig00000159,
      DI => blk00000003_sig0000015c,
      S => blk00000003_sig0000015a,
      O => blk00000003_sig00000155
    );
  blk00000003_blk00000113 : XORCY
    port map (
      CI => blk00000003_sig00000159,
      LI => blk00000003_sig0000015a,
      O => blk00000003_sig0000015b
    );
  blk00000003_blk00000112 : MUXCY
    port map (
      CI => blk00000003_sig00000146,
      DI => blk00000003_sig00000145,
      S => blk00000003_sig00000147,
      O => blk00000003_sig00000158
    );
  blk00000003_blk00000111 : MUXCY
    port map (
      CI => blk00000003_sig00000155,
      DI => blk00000003_sig00000140,
      S => blk00000003_sig00000156,
      O => blk00000003_sig00000152
    );
  blk00000003_blk00000110 : MUXCY
    port map (
      CI => blk00000003_sig00000152,
      DI => blk00000003_sig00000141,
      S => blk00000003_sig00000153,
      O => blk00000003_sig0000014f
    );
  blk00000003_blk0000010f : MUXCY
    port map (
      CI => blk00000003_sig0000014f,
      DI => blk00000003_sig00000142,
      S => blk00000003_sig00000150,
      O => blk00000003_sig0000014c
    );
  blk00000003_blk0000010e : MUXCY
    port map (
      CI => blk00000003_sig0000014c,
      DI => blk00000003_sig00000143,
      S => blk00000003_sig0000014d,
      O => blk00000003_sig00000149
    );
  blk00000003_blk0000010d : MUXCY
    port map (
      CI => blk00000003_sig00000149,
      DI => blk00000003_sig00000144,
      S => blk00000003_sig0000014a,
      O => blk00000003_sig00000146
    );
  blk00000003_blk0000010c : XORCY
    port map (
      CI => blk00000003_sig00000155,
      LI => blk00000003_sig00000156,
      O => blk00000003_sig00000157
    );
  blk00000003_blk0000010b : XORCY
    port map (
      CI => blk00000003_sig00000152,
      LI => blk00000003_sig00000153,
      O => blk00000003_sig00000154
    );
  blk00000003_blk0000010a : XORCY
    port map (
      CI => blk00000003_sig0000014f,
      LI => blk00000003_sig00000150,
      O => blk00000003_sig00000151
    );
  blk00000003_blk00000109 : XORCY
    port map (
      CI => blk00000003_sig0000014c,
      LI => blk00000003_sig0000014d,
      O => blk00000003_sig0000014e
    );
  blk00000003_blk00000108 : XORCY
    port map (
      CI => blk00000003_sig00000149,
      LI => blk00000003_sig0000014a,
      O => blk00000003_sig0000014b
    );
  blk00000003_blk00000107 : XORCY
    port map (
      CI => blk00000003_sig00000146,
      LI => blk00000003_sig00000147,
      O => blk00000003_sig00000148
    );
  blk00000003_blk00000106 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000012e,
      Q => blk00000003_sig0000006f
    );
  blk00000003_blk00000105 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000131,
      Q => blk00000003_sig00000145
    );
  blk00000003_blk00000104 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000134,
      Q => blk00000003_sig00000144
    );
  blk00000003_blk00000103 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000137,
      Q => blk00000003_sig00000143
    );
  blk00000003_blk00000102 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000013a,
      Q => blk00000003_sig00000142
    );
  blk00000003_blk00000101 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000013d,
      Q => blk00000003_sig00000141
    );
  blk00000003_blk00000100 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000013f,
      Q => blk00000003_sig00000140
    );
  blk00000003_blk000000ff : MUXCY
    port map (
      CI => NlwRenamedSig_OI_rfd,
      DI => blk00000003_sig00000121,
      S => blk00000003_sig0000013e,
      O => blk00000003_sig0000013b
    );
  blk00000003_blk000000fe : XORCY
    port map (
      CI => NlwRenamedSig_OI_rfd,
      LI => blk00000003_sig0000013e,
      O => blk00000003_sig0000013f
    );
  blk00000003_blk000000fd : MUXCY
    port map (
      CI => blk00000003_sig0000012d,
      DI => blk00000003_sig00000031,
      S => NlwRenamedSig_OI_rfd,
      O => NLW_blk00000003_blk000000fd_O_UNCONNECTED
    );
  blk00000003_blk000000fc : MUXCY
    port map (
      CI => blk00000003_sig0000013b,
      DI => blk00000003_sig00000031,
      S => blk00000003_sig0000013c,
      O => blk00000003_sig00000138
    );
  blk00000003_blk000000fb : MUXCY
    port map (
      CI => blk00000003_sig00000138,
      DI => blk00000003_sig00000031,
      S => blk00000003_sig00000139,
      O => blk00000003_sig00000135
    );
  blk00000003_blk000000fa : MUXCY
    port map (
      CI => blk00000003_sig00000135,
      DI => blk00000003_sig00000031,
      S => blk00000003_sig00000136,
      O => blk00000003_sig00000132
    );
  blk00000003_blk000000f9 : MUXCY
    port map (
      CI => blk00000003_sig00000132,
      DI => blk00000003_sig00000031,
      S => blk00000003_sig00000133,
      O => blk00000003_sig0000012f
    );
  blk00000003_blk000000f8 : MUXCY
    port map (
      CI => blk00000003_sig0000012f,
      DI => blk00000003_sig00000031,
      S => blk00000003_sig00000130,
      O => blk00000003_sig0000012d
    );
  blk00000003_blk000000f7 : XORCY
    port map (
      CI => blk00000003_sig0000013b,
      LI => blk00000003_sig0000013c,
      O => blk00000003_sig0000013d
    );
  blk00000003_blk000000f6 : XORCY
    port map (
      CI => blk00000003_sig00000138,
      LI => blk00000003_sig00000139,
      O => blk00000003_sig0000013a
    );
  blk00000003_blk000000f5 : XORCY
    port map (
      CI => blk00000003_sig00000135,
      LI => blk00000003_sig00000136,
      O => blk00000003_sig00000137
    );
  blk00000003_blk000000f4 : XORCY
    port map (
      CI => blk00000003_sig00000132,
      LI => blk00000003_sig00000133,
      O => blk00000003_sig00000134
    );
  blk00000003_blk000000f3 : XORCY
    port map (
      CI => blk00000003_sig0000012f,
      LI => blk00000003_sig00000130,
      O => blk00000003_sig00000131
    );
  blk00000003_blk000000f2 : XORCY
    port map (
      CI => blk00000003_sig0000012d,
      LI => NlwRenamedSig_OI_rfd,
      O => blk00000003_sig0000012e
    );
  blk00000003_blk000000f1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(0),
      Q => blk00000003_sig0000012c
    );
  blk00000003_blk000000f0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(1),
      Q => blk00000003_sig0000012b
    );
  blk00000003_blk000000ef : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(2),
      Q => blk00000003_sig0000012a
    );
  blk00000003_blk000000ee : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(3),
      Q => blk00000003_sig00000129
    );
  blk00000003_blk000000ed : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(4),
      Q => blk00000003_sig00000128
    );
  blk00000003_blk000000ec : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(5),
      Q => blk00000003_sig00000127
    );
  blk00000003_blk000000eb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(6),
      Q => blk00000003_sig00000126
    );
  blk00000003_blk000000ea : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(7),
      Q => blk00000003_sig00000125
    );
  blk00000003_blk000000e9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(8),
      Q => blk00000003_sig00000124
    );
  blk00000003_blk000000e8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(9),
      Q => blk00000003_sig00000123
    );
  blk00000003_blk000000e7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(10),
      Q => blk00000003_sig00000122
    );
  blk00000003_blk000000e6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(11),
      Q => blk00000003_sig00000121
    );
  blk00000003_blk000000e5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000011a,
      Q => blk00000003_sig00000120
    );
  blk00000003_blk000000e4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000119,
      Q => blk00000003_sig0000011f
    );
  blk00000003_blk000000e3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000118,
      Q => blk00000003_sig0000011e
    );
  blk00000003_blk000000e2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000117,
      Q => blk00000003_sig0000011d
    );
  blk00000003_blk000000e1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000116,
      Q => blk00000003_sig0000011c
    );
  blk00000003_blk000000e0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000115,
      Q => blk00000003_sig0000011b
    );
  blk00000003_blk000000df : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000114,
      Q => blk00000003_sig0000011a
    );
  blk00000003_blk000000de : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000113,
      Q => blk00000003_sig00000119
    );
  blk00000003_blk000000dd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000112,
      Q => blk00000003_sig00000118
    );
  blk00000003_blk000000dc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000111,
      Q => blk00000003_sig00000117
    );
  blk00000003_blk000000db : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000110,
      Q => blk00000003_sig00000116
    );
  blk00000003_blk000000da : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000010f,
      Q => blk00000003_sig00000115
    );
  blk00000003_blk000000d9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000010e,
      Q => blk00000003_sig00000114
    );
  blk00000003_blk000000d8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000010d,
      Q => blk00000003_sig00000113
    );
  blk00000003_blk000000d7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000010c,
      Q => blk00000003_sig00000112
    );
  blk00000003_blk000000d6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000010b,
      Q => blk00000003_sig00000111
    );
  blk00000003_blk000000d5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000010a,
      Q => blk00000003_sig00000110
    );
  blk00000003_blk000000d4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000109,
      Q => blk00000003_sig0000010f
    );
  blk00000003_blk000000d3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000108,
      Q => blk00000003_sig0000010e
    );
  blk00000003_blk000000d2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000107,
      Q => blk00000003_sig0000010d
    );
  blk00000003_blk000000d1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000106,
      Q => blk00000003_sig0000010c
    );
  blk00000003_blk000000d0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000105,
      Q => blk00000003_sig0000010b
    );
  blk00000003_blk000000cf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000104,
      Q => blk00000003_sig0000010a
    );
  blk00000003_blk000000ce : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000103,
      Q => blk00000003_sig00000109
    );
  blk00000003_blk000000cd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000102,
      Q => blk00000003_sig00000108
    );
  blk00000003_blk000000cc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000101,
      Q => blk00000003_sig00000107
    );
  blk00000003_blk000000cb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000100,
      Q => blk00000003_sig00000106
    );
  blk00000003_blk000000ca : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ff,
      Q => blk00000003_sig00000105
    );
  blk00000003_blk000000c9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000fe,
      Q => blk00000003_sig00000104
    );
  blk00000003_blk000000c8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000fd,
      Q => blk00000003_sig00000103
    );
  blk00000003_blk000000c7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000fc,
      Q => blk00000003_sig00000102
    );
  blk00000003_blk000000c6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000fb,
      Q => blk00000003_sig00000101
    );
  blk00000003_blk000000c5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000fa,
      Q => blk00000003_sig00000100
    );
  blk00000003_blk000000c4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f9,
      Q => blk00000003_sig000000ff
    );
  blk00000003_blk000000c3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f8,
      Q => blk00000003_sig000000fe
    );
  blk00000003_blk000000c2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f7,
      Q => blk00000003_sig000000fd
    );
  blk00000003_blk000000c1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f6,
      Q => blk00000003_sig000000fc
    );
  blk00000003_blk000000c0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f5,
      Q => blk00000003_sig000000fb
    );
  blk00000003_blk000000bf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f4,
      Q => blk00000003_sig000000fa
    );
  blk00000003_blk000000be : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f3,
      Q => blk00000003_sig000000f9
    );
  blk00000003_blk000000bd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f2,
      Q => blk00000003_sig000000f8
    );
  blk00000003_blk000000bc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f1,
      Q => blk00000003_sig000000f7
    );
  blk00000003_blk000000bb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f0,
      Q => blk00000003_sig000000f6
    );
  blk00000003_blk000000ba : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ef,
      Q => blk00000003_sig000000f5
    );
  blk00000003_blk000000b9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ee,
      Q => blk00000003_sig000000f4
    );
  blk00000003_blk000000b8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ed,
      Q => blk00000003_sig000000f3
    );
  blk00000003_blk000000b7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ec,
      Q => blk00000003_sig000000f2
    );
  blk00000003_blk000000b6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000eb,
      Q => blk00000003_sig000000f1
    );
  blk00000003_blk000000b5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ea,
      Q => blk00000003_sig000000f0
    );
  blk00000003_blk000000b4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e9,
      Q => blk00000003_sig000000ef
    );
  blk00000003_blk000000b3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e8,
      Q => blk00000003_sig000000ee
    );
  blk00000003_blk000000b2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e7,
      Q => blk00000003_sig000000ed
    );
  blk00000003_blk000000b1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e6,
      Q => blk00000003_sig000000ec
    );
  blk00000003_blk000000b0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e5,
      Q => blk00000003_sig000000eb
    );
  blk00000003_blk000000af : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e4,
      Q => blk00000003_sig000000ea
    );
  blk00000003_blk000000ae : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e3,
      Q => blk00000003_sig000000e9
    );
  blk00000003_blk000000ad : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e2,
      Q => blk00000003_sig000000e8
    );
  blk00000003_blk000000ac : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e1,
      Q => blk00000003_sig000000e7
    );
  blk00000003_blk000000ab : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e0,
      Q => blk00000003_sig000000e6
    );
  blk00000003_blk000000aa : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000df,
      Q => blk00000003_sig000000e5
    );
  blk00000003_blk000000a9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000de,
      Q => blk00000003_sig000000e4
    );
  blk00000003_blk000000a8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000dd,
      Q => blk00000003_sig000000e3
    );
  blk00000003_blk000000a7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000dc,
      Q => blk00000003_sig000000e2
    );
  blk00000003_blk000000a6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000db,
      Q => blk00000003_sig000000e1
    );
  blk00000003_blk000000a5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000da,
      Q => blk00000003_sig000000e0
    );
  blk00000003_blk000000a4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d9,
      Q => blk00000003_sig000000df
    );
  blk00000003_blk000000a3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d8,
      Q => blk00000003_sig000000de
    );
  blk00000003_blk000000a2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d7,
      Q => blk00000003_sig000000dd
    );
  blk00000003_blk000000a1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d6,
      Q => blk00000003_sig000000dc
    );
  blk00000003_blk000000a0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d5,
      Q => blk00000003_sig000000db
    );
  blk00000003_blk0000009f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d4,
      Q => blk00000003_sig000000da
    );
  blk00000003_blk0000009e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d3,
      Q => blk00000003_sig000000d9
    );
  blk00000003_blk0000009d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d2,
      Q => blk00000003_sig000000d8
    );
  blk00000003_blk0000009c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d1,
      Q => blk00000003_sig000000d7
    );
  blk00000003_blk0000009b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d0,
      Q => blk00000003_sig000000d6
    );
  blk00000003_blk0000009a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000cf,
      Q => blk00000003_sig000000d5
    );
  blk00000003_blk00000099 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ce,
      Q => blk00000003_sig000000d4
    );
  blk00000003_blk00000098 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000cd,
      Q => blk00000003_sig000000d3
    );
  blk00000003_blk00000097 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000cc,
      Q => blk00000003_sig000000d2
    );
  blk00000003_blk00000096 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000cb,
      Q => blk00000003_sig000000d1
    );
  blk00000003_blk00000095 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ca,
      Q => blk00000003_sig000000d0
    );
  blk00000003_blk00000094 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c9,
      Q => blk00000003_sig000000cf
    );
  blk00000003_blk00000093 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c8,
      Q => blk00000003_sig000000ce
    );
  blk00000003_blk00000092 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c7,
      Q => blk00000003_sig000000cd
    );
  blk00000003_blk00000091 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c6,
      Q => blk00000003_sig000000cc
    );
  blk00000003_blk00000090 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c5,
      Q => blk00000003_sig000000cb
    );
  blk00000003_blk0000008f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c4,
      Q => blk00000003_sig000000ca
    );
  blk00000003_blk0000008e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c3,
      Q => blk00000003_sig000000c9
    );
  blk00000003_blk0000008d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c2,
      Q => blk00000003_sig000000c8
    );
  blk00000003_blk0000008c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c1,
      Q => blk00000003_sig000000c7
    );
  blk00000003_blk0000008b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c0,
      Q => blk00000003_sig000000c6
    );
  blk00000003_blk0000008a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000bf,
      Q => blk00000003_sig000000c5
    );
  blk00000003_blk00000089 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000be,
      Q => blk00000003_sig000000c4
    );
  blk00000003_blk00000088 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000bd,
      Q => blk00000003_sig000000c3
    );
  blk00000003_blk00000087 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000bc,
      Q => blk00000003_sig000000c2
    );
  blk00000003_blk00000086 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000bb,
      Q => blk00000003_sig000000c1
    );
  blk00000003_blk00000085 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ba,
      Q => blk00000003_sig000000c0
    );
  blk00000003_blk00000084 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b9,
      Q => blk00000003_sig000000bf
    );
  blk00000003_blk00000083 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b8,
      Q => blk00000003_sig000000be
    );
  blk00000003_blk00000082 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b7,
      Q => blk00000003_sig000000bd
    );
  blk00000003_blk00000081 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b6,
      Q => blk00000003_sig000000bc
    );
  blk00000003_blk00000080 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b5,
      Q => blk00000003_sig000000bb
    );
  blk00000003_blk0000007f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b4,
      Q => blk00000003_sig000000ba
    );
  blk00000003_blk0000007e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b3,
      Q => blk00000003_sig000000b9
    );
  blk00000003_blk0000007d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b2,
      Q => blk00000003_sig000000b8
    );
  blk00000003_blk0000007c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b1,
      Q => blk00000003_sig000000b7
    );
  blk00000003_blk0000007b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b0,
      Q => blk00000003_sig000000b6
    );
  blk00000003_blk0000007a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000af,
      Q => blk00000003_sig000000b5
    );
  blk00000003_blk00000079 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ae,
      Q => blk00000003_sig000000b4
    );
  blk00000003_blk00000078 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ad,
      Q => blk00000003_sig000000b3
    );
  blk00000003_blk00000077 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ac,
      Q => blk00000003_sig000000b2
    );
  blk00000003_blk00000076 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ab,
      Q => blk00000003_sig000000b1
    );
  blk00000003_blk00000075 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000aa,
      Q => blk00000003_sig000000b0
    );
  blk00000003_blk00000074 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a9,
      Q => blk00000003_sig000000af
    );
  blk00000003_blk00000073 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a8,
      Q => blk00000003_sig000000ae
    );
  blk00000003_blk00000072 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a7,
      Q => blk00000003_sig000000ad
    );
  blk00000003_blk00000071 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a6,
      Q => blk00000003_sig000000ac
    );
  blk00000003_blk00000070 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a5,
      Q => blk00000003_sig000000ab
    );
  blk00000003_blk0000006f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a4,
      Q => blk00000003_sig000000aa
    );
  blk00000003_blk0000006e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a3,
      Q => blk00000003_sig000000a9
    );
  blk00000003_blk0000006d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a2,
      Q => blk00000003_sig000000a8
    );
  blk00000003_blk0000006c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a1,
      Q => blk00000003_sig000000a7
    );
  blk00000003_blk0000006b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a0,
      Q => blk00000003_sig000000a6
    );
  blk00000003_blk0000006a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000009f,
      Q => blk00000003_sig000000a5
    );
  blk00000003_blk00000069 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000009e,
      Q => blk00000003_sig000000a4
    );
  blk00000003_blk00000068 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000009d,
      Q => blk00000003_sig000000a3
    );
  blk00000003_blk00000067 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000009c,
      Q => blk00000003_sig000000a2
    );
  blk00000003_blk00000066 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000009b,
      Q => blk00000003_sig000000a1
    );
  blk00000003_blk00000065 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000009a,
      Q => blk00000003_sig000000a0
    );
  blk00000003_blk00000064 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000099,
      Q => blk00000003_sig0000009f
    );
  blk00000003_blk00000063 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000098,
      Q => blk00000003_sig0000009e
    );
  blk00000003_blk00000062 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000097,
      Q => blk00000003_sig0000009d
    );
  blk00000003_blk00000061 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000096,
      Q => blk00000003_sig0000009c
    );
  blk00000003_blk00000060 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000095,
      Q => blk00000003_sig0000009b
    );
  blk00000003_blk0000005f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000094,
      Q => blk00000003_sig0000009a
    );
  blk00000003_blk0000005e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000093,
      Q => blk00000003_sig00000099
    );
  blk00000003_blk0000005d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000092,
      Q => blk00000003_sig00000098
    );
  blk00000003_blk0000005c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000091,
      Q => blk00000003_sig00000097
    );
  blk00000003_blk0000005b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000090,
      Q => blk00000003_sig00000096
    );
  blk00000003_blk0000005a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000008f,
      Q => blk00000003_sig00000095
    );
  blk00000003_blk00000059 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000008e,
      Q => blk00000003_sig00000094
    );
  blk00000003_blk00000058 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000008d,
      Q => blk00000003_sig00000093
    );
  blk00000003_blk00000057 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000008c,
      Q => blk00000003_sig00000092
    );
  blk00000003_blk00000056 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000008b,
      Q => blk00000003_sig00000091
    );
  blk00000003_blk00000055 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000008a,
      Q => blk00000003_sig00000090
    );
  blk00000003_blk00000054 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000089,
      Q => blk00000003_sig0000008f
    );
  blk00000003_blk00000053 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000088,
      Q => blk00000003_sig0000008e
    );
  blk00000003_blk00000052 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000087,
      Q => blk00000003_sig0000008d
    );
  blk00000003_blk00000051 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000086,
      Q => blk00000003_sig0000008c
    );
  blk00000003_blk00000050 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000085,
      Q => blk00000003_sig0000008b
    );
  blk00000003_blk0000004f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000084,
      Q => blk00000003_sig0000008a
    );
  blk00000003_blk0000004e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000083,
      Q => blk00000003_sig00000089
    );
  blk00000003_blk0000004d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000082,
      Q => blk00000003_sig00000088
    );
  blk00000003_blk0000004c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000081,
      Q => blk00000003_sig00000087
    );
  blk00000003_blk0000004b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000080,
      Q => blk00000003_sig00000086
    );
  blk00000003_blk0000004a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007f,
      Q => blk00000003_sig00000085
    );
  blk00000003_blk00000049 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007e,
      Q => blk00000003_sig00000084
    );
  blk00000003_blk00000048 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007d,
      Q => blk00000003_sig00000083
    );
  blk00000003_blk00000047 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007c,
      Q => blk00000003_sig00000082
    );
  blk00000003_blk00000046 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007b,
      Q => blk00000003_sig00000081
    );
  blk00000003_blk00000045 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007a,
      Q => blk00000003_sig00000080
    );
  blk00000003_blk00000044 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000079,
      Q => blk00000003_sig0000007f
    );
  blk00000003_blk00000043 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(5),
      Q => blk00000003_sig0000007e
    );
  blk00000003_blk00000042 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(4),
      Q => blk00000003_sig0000007d
    );
  blk00000003_blk00000041 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(3),
      Q => blk00000003_sig0000007c
    );
  blk00000003_blk00000040 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(2),
      Q => blk00000003_sig0000007b
    );
  blk00000003_blk0000003f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(1),
      Q => blk00000003_sig0000007a
    );
  blk00000003_blk0000003e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(0),
      Q => blk00000003_sig00000079
    );
  blk00000003_blk0000003d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000034,
      Q => blk00000003_sig00000078
    );
  blk00000003_blk0000003c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000051,
      Q => blk00000003_sig00000077
    );
  blk00000003_blk0000003b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000004f,
      Q => blk00000003_sig00000076
    );
  blk00000003_blk0000003a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000004d,
      Q => blk00000003_sig00000075
    );
  blk00000003_blk00000039 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000004b,
      Q => blk00000003_sig00000074
    );
  blk00000003_blk00000038 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000049,
      Q => blk00000003_sig00000073
    );
  blk00000003_blk00000037 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000047,
      Q => blk00000003_sig00000072
    );
  blk00000003_blk00000036 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000070,
      Q => blk00000003_sig00000071
    );
  blk00000003_blk00000035 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006f,
      Q => blk00000003_sig0000006e
    );
  blk00000003_blk00000034 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006e,
      Q => blk00000003_sig0000006c
    );
  blk00000003_blk00000033 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006d,
      Q => blk00000003_sig0000006b
    );
  blk00000003_blk00000032 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006c,
      Q => blk00000003_sig00000069
    );
  blk00000003_blk00000031 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006b,
      Q => blk00000003_sig00000068
    );
  blk00000003_blk00000030 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006a,
      Q => blk00000003_sig00000067
    );
  blk00000003_blk0000002f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000069,
      Q => blk00000003_sig0000005d
    );
  blk00000003_blk0000002e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000068,
      Q => blk00000003_sig0000005c
    );
  blk00000003_blk0000002d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000067,
      Q => blk00000003_sig0000005b
    );
  blk00000003_blk0000002c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000066,
      Q => blk00000003_sig0000005a
    );
  blk00000003_blk0000002b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000064,
      Q => blk00000003_sig00000065
    );
  blk00000003_blk0000002a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000063,
      Q => blk00000003_sig00000057
    );
  blk00000003_blk00000029 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000062,
      Q => blk00000003_sig00000056
    );
  blk00000003_blk00000028 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000061,
      Q => blk00000003_sig00000055
    );
  blk00000003_blk00000027 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000060,
      Q => blk00000003_sig00000054
    );
  blk00000003_blk00000026 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000005f,
      Q => blk00000003_sig00000053
    );
  blk00000003_blk00000025 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000005e,
      Q => blk00000003_sig00000052
    );
  blk00000003_blk00000024 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000005d,
      Q => blk00000003_sig00000050
    );
  blk00000003_blk00000023 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000005c,
      Q => blk00000003_sig0000004e
    );
  blk00000003_blk00000022 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000005b,
      Q => blk00000003_sig0000004c
    );
  blk00000003_blk00000021 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000005a,
      Q => blk00000003_sig0000004a
    );
  blk00000003_blk00000020 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000059,
      Q => blk00000003_sig00000048
    );
  blk00000003_blk0000001f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000057,
      Q => blk00000003_sig00000058
    );
  blk00000003_blk0000001e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000056,
      Q => blk00000003_sig00000044
    );
  blk00000003_blk0000001d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000055,
      Q => blk00000003_sig00000043
    );
  blk00000003_blk0000001c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000054,
      Q => blk00000003_sig00000042
    );
  blk00000003_blk0000001b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000053,
      Q => blk00000003_sig00000041
    );
  blk00000003_blk0000001a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000052,
      Q => blk00000003_sig00000040
    );
  blk00000003_blk00000019 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000050,
      Q => blk00000003_sig00000051
    );
  blk00000003_blk00000018 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000004e,
      Q => blk00000003_sig0000004f
    );
  blk00000003_blk00000017 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000004c,
      Q => blk00000003_sig0000004d
    );
  blk00000003_blk00000016 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000004a,
      Q => blk00000003_sig0000004b
    );
  blk00000003_blk00000015 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000048,
      Q => blk00000003_sig00000049
    );
  blk00000003_blk00000014 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000046,
      Q => blk00000003_sig00000047
    );
  blk00000003_blk00000013 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000044,
      Q => blk00000003_sig00000045
    );
  blk00000003_blk00000012 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000043,
      Q => blk00000003_sig0000003e
    );
  blk00000003_blk00000011 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000042,
      Q => blk00000003_sig0000003d
    );
  blk00000003_blk00000010 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000041,
      Q => blk00000003_sig0000003c
    );
  blk00000003_blk0000000f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000040,
      Q => blk00000003_sig0000003b
    );
  blk00000003_blk0000000e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000003e,
      Q => blk00000003_sig0000003f
    );
  blk00000003_blk0000000d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000003d,
      Q => blk00000003_sig00000039
    );
  blk00000003_blk0000000c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000003c,
      Q => blk00000003_sig00000038
    );
  blk00000003_blk0000000b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000003b,
      Q => blk00000003_sig00000037
    );
  blk00000003_blk0000000a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000039,
      Q => blk00000003_sig0000003a
    );
  blk00000003_blk00000009 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000038,
      Q => blk00000003_sig00000035
    );
  blk00000003_blk00000008 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000037,
      Q => blk00000003_sig00000033
    );
  blk00000003_blk00000007 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000035,
      Q => blk00000003_sig00000036
    );
  blk00000003_blk00000006 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000033,
      Q => blk00000003_sig00000034
    );
  blk00000003_blk00000005 : VCC
    port map (
      P => NlwRenamedSig_OI_rfd
    );
  blk00000003_blk00000004 : GND
    port map (
      G => blk00000003_sig00000031
    );

end STRUCTURE;

-- synthesis translate_on

-------------------------------------------------------------------
-- System Generator version 13.2 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
package conv_pkg is
    constant simulating : boolean := false
      -- synopsys translate_off
        or true
      -- synopsys translate_on
    ;
    constant xlUnsigned : integer := 1;
    constant xlSigned : integer := 2;
    constant xlWrap : integer := 1;
    constant xlSaturate : integer := 2;
    constant xlTruncate : integer := 1;
    constant xlRound : integer := 2;
    constant xlRoundBanker : integer := 3;
    constant xlAddMode : integer := 1;
    constant xlSubMode : integer := 2;
    attribute black_box : boolean;
    attribute syn_black_box : boolean;
    attribute fpga_dont_touch: string;
    attribute box_type :  string;
    attribute keep : string;
    attribute syn_keep : boolean;
    function std_logic_vector_to_unsigned(inp : std_logic_vector) return unsigned;
    function unsigned_to_std_logic_vector(inp : unsigned) return std_logic_vector;
    function std_logic_vector_to_signed(inp : std_logic_vector) return signed;
    function signed_to_std_logic_vector(inp : signed) return std_logic_vector;
    function unsigned_to_signed(inp : unsigned) return signed;
    function signed_to_unsigned(inp : signed) return unsigned;
    function pos(inp : std_logic_vector; arith : INTEGER) return boolean;
    function all_same(inp: std_logic_vector) return boolean;
    function all_zeros(inp: std_logic_vector) return boolean;
    function is_point_five(inp: std_logic_vector) return boolean;
    function all_ones(inp: std_logic_vector) return boolean;
    function convert_type (inp : std_logic_vector; old_width, old_bin_pt,
                           old_arith, new_width, new_bin_pt, new_arith,
                           quantization, overflow : INTEGER)
        return std_logic_vector;
    function cast (inp : std_logic_vector; old_bin_pt,
                   new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector;
    function vec_slice (inp : std_logic_vector; upper, lower : INTEGER)
        return std_logic_vector;
    function s2u_slice (inp : signed; upper, lower : INTEGER)
        return unsigned;
    function u2u_slice (inp : unsigned; upper, lower : INTEGER)
        return unsigned;
    function s2s_cast (inp : signed; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return signed;
    function u2s_cast (inp : unsigned; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return signed;
    function s2u_cast (inp : signed; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return unsigned;
    function u2u_cast (inp : unsigned; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return unsigned;
    function u2v_cast (inp : unsigned; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return std_logic_vector;
    function s2v_cast (inp : signed; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return std_logic_vector;
    function trunc (inp : std_logic_vector; old_width, old_bin_pt, old_arith,
                    new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector;
    function round_towards_inf (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt,
                                new_arith : INTEGER) return std_logic_vector;
    function round_towards_even (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt,
                                new_arith : INTEGER) return std_logic_vector;
    function max_signed(width : INTEGER) return std_logic_vector;
    function min_signed(width : INTEGER) return std_logic_vector;
    function saturation_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                              old_arith, new_width, new_bin_pt, new_arith
                              : INTEGER) return std_logic_vector;
    function wrap_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                        old_arith, new_width, new_bin_pt, new_arith : INTEGER)
                        return std_logic_vector;
    function fractional_bits(a_bin_pt, b_bin_pt: INTEGER) return INTEGER;
    function integer_bits(a_width, a_bin_pt, b_width, b_bin_pt: INTEGER)
        return INTEGER;
    function sign_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector;
    function zero_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector;
    function zero_ext(inp : std_logic; new_width : INTEGER)
        return std_logic_vector;
    function extend_MSB(inp : std_logic_vector; new_width, arith : INTEGER)
        return std_logic_vector;
    function align_input(inp : std_logic_vector; old_width, delta, new_arith,
                          new_width: INTEGER)
        return std_logic_vector;
    function pad_LSB(inp : std_logic_vector; new_width: integer)
        return std_logic_vector;
    function pad_LSB(inp : std_logic_vector; new_width, arith : integer)
        return std_logic_vector;
    function max(L, R: INTEGER) return INTEGER;
    function min(L, R: INTEGER) return INTEGER;
    function "="(left,right: STRING) return boolean;
    function boolean_to_signed (inp : boolean; width: integer)
        return signed;
    function boolean_to_unsigned (inp : boolean; width: integer)
        return unsigned;
    function boolean_to_vector (inp : boolean)
        return std_logic_vector;
    function std_logic_to_vector (inp : std_logic)
        return std_logic_vector;
    function integer_to_std_logic_vector (inp : integer;  width, arith : integer)
        return std_logic_vector;
    function std_logic_vector_to_integer (inp : std_logic_vector;  arith : integer)
        return integer;
    function std_logic_to_integer(constant inp : std_logic := '0')
        return integer;
    function bin_string_element_to_std_logic_vector (inp : string;  width, index : integer)
        return std_logic_vector;
    function bin_string_to_std_logic_vector (inp : string)
        return std_logic_vector;
    function hex_string_to_std_logic_vector (inp : string; width : integer)
        return std_logic_vector;
    function makeZeroBinStr (width : integer) return STRING;
    function and_reduce(inp: std_logic_vector) return std_logic;
    -- synopsys translate_off
    function is_binary_string_invalid (inp : string)
        return boolean;
    function is_binary_string_undefined (inp : string)
        return boolean;
    function is_XorU(inp : std_logic_vector)
        return boolean;
    function to_real(inp : std_logic_vector; bin_pt : integer; arith : integer)
        return real;
    function std_logic_to_real(inp : std_logic; bin_pt : integer; arith : integer)
        return real;
    function real_to_std_logic_vector (inp : real;  width, bin_pt, arith : integer)
        return std_logic_vector;
    function real_string_to_std_logic_vector (inp : string;  width, bin_pt, arith : integer)
        return std_logic_vector;
    constant display_precision : integer := 20;
    function real_to_string (inp : real) return string;
    function valid_bin_string(inp : string) return boolean;
    function std_logic_vector_to_bin_string(inp : std_logic_vector) return string;
    function std_logic_to_bin_string(inp : std_logic) return string;
    function std_logic_vector_to_bin_string_w_point(inp : std_logic_vector; bin_pt : integer)
        return string;
    function real_to_bin_string(inp : real;  width, bin_pt, arith : integer)
        return string;
    type stdlogic_to_char_t is array(std_logic) of character;
    constant to_char : stdlogic_to_char_t := (
        'U' => 'U',
        'X' => 'X',
        '0' => '0',
        '1' => '1',
        'Z' => 'Z',
        'W' => 'W',
        'L' => 'L',
        'H' => 'H',
        '-' => '-');
    -- synopsys translate_on
end conv_pkg;
package body conv_pkg is
    function std_logic_vector_to_unsigned(inp : std_logic_vector)
        return unsigned
    is
    begin
        return unsigned (inp);
    end;
    function unsigned_to_std_logic_vector(inp : unsigned)
        return std_logic_vector
    is
    begin
        return std_logic_vector(inp);
    end;
    function std_logic_vector_to_signed(inp : std_logic_vector)
        return signed
    is
    begin
        return  signed (inp);
    end;
    function signed_to_std_logic_vector(inp : signed)
        return std_logic_vector
    is
    begin
        return std_logic_vector(inp);
    end;
    function unsigned_to_signed (inp : unsigned)
        return signed
    is
    begin
        return signed(std_logic_vector(inp));
    end;
    function signed_to_unsigned (inp : signed)
        return unsigned
    is
    begin
        return unsigned(std_logic_vector(inp));
    end;
    function pos(inp : std_logic_vector; arith : INTEGER)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        if arith = xlUnsigned then
            return true;
        else
            if vec(width-1) = '0' then
                return true;
            else
                return false;
            end if;
        end if;
        return true;
    end;
    function max_signed(width : INTEGER)
        return std_logic_vector
    is
        variable ones : std_logic_vector(width-2 downto 0);
        variable result : std_logic_vector(width-1 downto 0);
    begin
        ones := (others => '1');
        result(width-1) := '0';
        result(width-2 downto 0) := ones;
        return result;
    end;
    function min_signed(width : INTEGER)
        return std_logic_vector
    is
        variable zeros : std_logic_vector(width-2 downto 0);
        variable result : std_logic_vector(width-1 downto 0);
    begin
        zeros := (others => '0');
        result(width-1) := '1';
        result(width-2 downto 0) := zeros;
        return result;
    end;
    function and_reduce(inp: std_logic_vector) return std_logic
    is
        variable result: std_logic;
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        result := vec(0);
        if width > 1 then
            for i in 1 to width-1 loop
                result := result and vec(i);
            end loop;
        end if;
        return result;
    end;
    function all_same(inp: std_logic_vector) return boolean
    is
        variable result: boolean;
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        result := true;
        if width > 0 then
            for i in 1 to width-1 loop
                if vec(i) /= vec(0) then
                    result := false;
                end if;
            end loop;
        end if;
        return result;
    end;
    function all_zeros(inp: std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable zero : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        zero := (others => '0');
        vec := inp;
        -- synopsys translate_off
        if (is_XorU(vec)) then
            return false;
        end if;
         -- synopsys translate_on
        if (std_logic_vector_to_unsigned(vec) = std_logic_vector_to_unsigned(zero)) then
            result := true;
        else
            result := false;
        end if;
        return result;
    end;
    function is_point_five(inp: std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        vec := inp;
        -- synopsys translate_off
        if (is_XorU(vec)) then
            return false;
        end if;
         -- synopsys translate_on
        if (width > 1) then
           if ((vec(width-1) = '1') and (all_zeros(vec(width-2 downto 0)) = true)) then
               result := true;
           else
               result := false;
           end if;
        else
           if (vec(width-1) = '1') then
               result := true;
           else
               result := false;
           end if;
        end if;
        return result;
    end;
    function all_ones(inp: std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable one : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        one := (others => '1');
        vec := inp;
        -- synopsys translate_off
        if (is_XorU(vec)) then
            return false;
        end if;
         -- synopsys translate_on
        if (std_logic_vector_to_unsigned(vec) = std_logic_vector_to_unsigned(one)) then
            result := true;
        else
            result := false;
        end if;
        return result;
    end;
    function full_precision_num_width(quantization, overflow, old_width,
                                      old_bin_pt, old_arith,
                                      new_width, new_bin_pt, new_arith : INTEGER)
        return integer
    is
        variable result : integer;
    begin
        result := old_width + 2;
        return result;
    end;
    function quantized_num_width(quantization, overflow, old_width, old_bin_pt,
                                 old_arith, new_width, new_bin_pt, new_arith
                                 : INTEGER)
        return integer
    is
        variable right_of_dp, left_of_dp, result : integer;
    begin
        right_of_dp := max(new_bin_pt, old_bin_pt);
        left_of_dp := max((new_width - new_bin_pt), (old_width - old_bin_pt));
        result := (old_width + 2) + (new_bin_pt - old_bin_pt);
        return result;
    end;
    function convert_type (inp : std_logic_vector; old_width, old_bin_pt,
                           old_arith, new_width, new_bin_pt, new_arith,
                           quantization, overflow : INTEGER)
        return std_logic_vector
    is
        constant fp_width : integer :=
            full_precision_num_width(quantization, overflow, old_width,
                                     old_bin_pt, old_arith, new_width,
                                     new_bin_pt, new_arith);
        constant fp_bin_pt : integer := old_bin_pt;
        constant fp_arith : integer := old_arith;
        variable full_precision_result : std_logic_vector(fp_width-1 downto 0);
        constant q_width : integer :=
            quantized_num_width(quantization, overflow, old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt, new_arith);
        constant q_bin_pt : integer := new_bin_pt;
        constant q_arith : integer := old_arith;
        variable quantized_result : std_logic_vector(q_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        result := (others => '0');
        full_precision_result := cast(inp, old_bin_pt, fp_width, fp_bin_pt,
                                      fp_arith);
        if (quantization = xlRound) then
            quantized_result := round_towards_inf(full_precision_result,
                                                  fp_width, fp_bin_pt,
                                                  fp_arith, q_width, q_bin_pt,
                                                  q_arith);
        elsif (quantization = xlRoundBanker) then
            quantized_result := round_towards_even(full_precision_result,
                                                  fp_width, fp_bin_pt,
                                                  fp_arith, q_width, q_bin_pt,
                                                  q_arith);
        else
            quantized_result := trunc(full_precision_result, fp_width, fp_bin_pt,
                                      fp_arith, q_width, q_bin_pt, q_arith);
        end if;
        if (overflow = xlSaturate) then
            result := saturation_arith(quantized_result, q_width, q_bin_pt,
                                       q_arith, new_width, new_bin_pt, new_arith);
        else
             result := wrap_arith(quantized_result, q_width, q_bin_pt, q_arith,
                                  new_width, new_bin_pt, new_arith);
        end if;
        return result;
    end;
    function cast (inp : std_logic_vector; old_bin_pt, new_width,
                   new_bin_pt, new_arith : INTEGER)
        return std_logic_vector
    is
        constant old_width : integer := inp'length;
        constant left_of_dp : integer := (new_width - new_bin_pt)
                                         - (old_width - old_bin_pt);
        constant right_of_dp : integer := (new_bin_pt - old_bin_pt);
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable j   : integer;
    begin
        vec := inp;
        for i in new_width-1 downto 0 loop
            j := i - right_of_dp;
            if ( j > old_width-1) then
                if (new_arith = xlUnsigned) then
                    result(i) := '0';
                else
                    result(i) := vec(old_width-1);
                end if;
            elsif ( j >= 0) then
                result(i) := vec(j);
            else
                result(i) := '0';
            end if;
        end loop;
        return result;
    end;
    function vec_slice (inp : std_logic_vector; upper, lower : INTEGER)
      return std_logic_vector
    is
    begin
        return inp(upper downto lower);
    end;
    function s2u_slice (inp : signed; upper, lower : INTEGER)
      return unsigned
    is
    begin
        return unsigned(vec_slice(std_logic_vector(inp), upper, lower));
    end;
    function u2u_slice (inp : unsigned; upper, lower : INTEGER)
      return unsigned
    is
    begin
        return unsigned(vec_slice(std_logic_vector(inp), upper, lower));
    end;
    function s2s_cast (inp : signed; old_bin_pt, new_width, new_bin_pt : INTEGER)
        return signed
    is
    begin
        return signed(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlSigned));
    end;
    function s2u_cast (inp : signed; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return unsigned
    is
    begin
        return unsigned(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlSigned));
    end;
    function u2s_cast (inp : unsigned; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return signed
    is
    begin
        return signed(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlUnsigned));
    end;
    function u2u_cast (inp : unsigned; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return unsigned
    is
    begin
        return unsigned(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlUnsigned));
    end;
    function u2v_cast (inp : unsigned; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return std_logic_vector
    is
    begin
        return cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlUnsigned);
    end;
    function s2v_cast (inp : signed; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return std_logic_vector
    is
    begin
        return cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlSigned);
    end;
    function boolean_to_signed (inp : boolean; width : integer)
        return signed
    is
        variable result : signed(width - 1 downto 0);
    begin
        result := (others => '0');
        if inp then
          result(0) := '1';
        else
          result(0) := '0';
        end if;
        return result;
    end;
    function boolean_to_unsigned (inp : boolean; width : integer)
        return unsigned
    is
        variable result : unsigned(width - 1 downto 0);
    begin
        result := (others => '0');
        if inp then
          result(0) := '1';
        else
          result(0) := '0';
        end if;
        return result;
    end;
    function boolean_to_vector (inp : boolean)
        return std_logic_vector
    is
        variable result : std_logic_vector(1 - 1 downto 0);
    begin
        result := (others => '0');
        if inp then
          result(0) := '1';
        else
          result(0) := '0';
        end if;
        return result;
    end;
    function std_logic_to_vector (inp : std_logic)
        return std_logic_vector
    is
        variable result : std_logic_vector(1 - 1 downto 0);
    begin
        result(0) := inp;
        return result;
    end;
    function trunc (inp : std_logic_vector; old_width, old_bin_pt, old_arith,
                                new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector
    is
        constant right_of_dp : integer := (old_bin_pt - new_bin_pt);
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if right_of_dp >= 0 then
            if new_arith = xlUnsigned then
                result := zero_ext(vec(old_width-1 downto right_of_dp), new_width);
            else
                result := sign_ext(vec(old_width-1 downto right_of_dp), new_width);
            end if;
        else
            if new_arith = xlUnsigned then
                result := zero_ext(pad_LSB(vec, old_width +
                                           abs(right_of_dp)), new_width);
            else
                result := sign_ext(pad_LSB(vec, old_width +
                                           abs(right_of_dp)), new_width);
            end if;
        end if;
        return result;
    end;
    function round_towards_inf (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt, new_arith
                                : INTEGER)
        return std_logic_vector
    is
        constant right_of_dp : integer := (old_bin_pt - new_bin_pt);
        constant expected_new_width : integer :=  old_width - right_of_dp  + 1;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable one_or_zero : std_logic_vector(new_width-1 downto 0);
        variable truncated_val : std_logic_vector(new_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if right_of_dp >= 0 then
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            else
                truncated_val := sign_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            end if;
        else
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            else
                truncated_val := sign_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            end if;
        end if;
        one_or_zero := (others => '0');
        if (new_arith = xlSigned) then
            if (vec(old_width-1) = '0') then
                one_or_zero(0) := '1';
            end if;
            if (right_of_dp >= 2) and (right_of_dp <= old_width) then
                if (all_zeros(vec(right_of_dp-2 downto 0)) = false) then
                    one_or_zero(0) := '1';
                end if;
            end if;
            if (right_of_dp >= 1) and (right_of_dp <= old_width) then
                if vec(right_of_dp-1) = '0' then
                    one_or_zero(0) := '0';
                end if;
            else
                one_or_zero(0) := '0';
            end if;
        else
            if (right_of_dp >= 1) and (right_of_dp <= old_width) then
                one_or_zero(0) :=  vec(right_of_dp-1);
            end if;
        end if;
        if new_arith = xlSigned then
            result := signed_to_std_logic_vector(std_logic_vector_to_signed(truncated_val) +
                                                 std_logic_vector_to_signed(one_or_zero));
        else
            result := unsigned_to_std_logic_vector(std_logic_vector_to_unsigned(truncated_val) +
                                                  std_logic_vector_to_unsigned(one_or_zero));
        end if;
        return result;
    end;
    function round_towards_even (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt, new_arith
                                : INTEGER)
        return std_logic_vector
    is
        constant right_of_dp : integer := (old_bin_pt - new_bin_pt);
        constant expected_new_width : integer :=  old_width - right_of_dp  + 1;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable one_or_zero : std_logic_vector(new_width-1 downto 0);
        variable truncated_val : std_logic_vector(new_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if right_of_dp >= 0 then
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            else
                truncated_val := sign_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            end if;
        else
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            else
                truncated_val := sign_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            end if;
        end if;
        one_or_zero := (others => '0');
        if (right_of_dp >= 1) and (right_of_dp <= old_width) then
            if (is_point_five(vec(right_of_dp-1 downto 0)) = false) then
                one_or_zero(0) :=  vec(right_of_dp-1);
            else
                one_or_zero(0) :=  vec(right_of_dp);
            end if;
        end if;
        if new_arith = xlSigned then
            result := signed_to_std_logic_vector(std_logic_vector_to_signed(truncated_val) +
                                                 std_logic_vector_to_signed(one_or_zero));
        else
            result := unsigned_to_std_logic_vector(std_logic_vector_to_unsigned(truncated_val) +
                                                  std_logic_vector_to_unsigned(one_or_zero));
        end if;
        return result;
    end;
    function saturation_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                              old_arith, new_width, new_bin_pt, new_arith
                              : INTEGER)
        return std_logic_vector
    is
        constant left_of_dp : integer := (old_width - old_bin_pt) -
                                         (new_width - new_bin_pt);
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable overflow : boolean;
    begin
        vec := inp;
        overflow := true;
        result := (others => '0');
        if (new_width >= old_width) then
            overflow := false;
        end if;
        if ((old_arith = xlSigned and new_arith = xlSigned) and (old_width > new_width)) then
            if all_same(vec(old_width-1 downto new_width-1)) then
                overflow := false;
            end if;
        end if;
        if (old_arith = xlSigned and new_arith = xlUnsigned) then
            if (old_width > new_width) then
                if all_zeros(vec(old_width-1 downto new_width)) then
                    overflow := false;
                end if;
            else
                if (old_width = new_width) then
                    if (vec(new_width-1) = '0') then
                        overflow := false;
                    end if;
                end if;
            end if;
        end if;
        if (old_arith = xlUnsigned and new_arith = xlUnsigned) then
            if (old_width > new_width) then
                if all_zeros(vec(old_width-1 downto new_width)) then
                    overflow := false;
                end if;
            else
                if (old_width = new_width) then
                    overflow := false;
                end if;
            end if;
        end if;
        if ((old_arith = xlUnsigned and new_arith = xlSigned) and (old_width > new_width)) then
            if all_same(vec(old_width-1 downto new_width-1)) then
                overflow := false;
            end if;
        end if;
        if overflow then
            if new_arith = xlSigned then
                if vec(old_width-1) = '0' then
                    result := max_signed(new_width);
                else
                    result := min_signed(new_width);
                end if;
            else
                if ((old_arith = xlSigned) and vec(old_width-1) = '1') then
                    result := (others => '0');
                else
                    result := (others => '1');
                end if;
            end if;
        else
            if (old_arith = xlSigned) and (new_arith = xlUnsigned) then
                if (vec(old_width-1) = '1') then
                    vec := (others => '0');
                end if;
            end if;
            if new_width <= old_width then
                result := vec(new_width-1 downto 0);
            else
                if new_arith = xlUnsigned then
                    result := zero_ext(vec, new_width);
                else
                    result := sign_ext(vec, new_width);
                end if;
            end if;
        end if;
        return result;
    end;
   function wrap_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                       old_arith, new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector
    is
        variable result : std_logic_vector(new_width-1 downto 0);
        variable result_arith : integer;
    begin
        if (old_arith = xlSigned) and (new_arith = xlUnsigned) then
            result_arith := xlSigned;
        end if;
        result := cast(inp, old_bin_pt, new_width, new_bin_pt, result_arith);
        return result;
    end;
    function fractional_bits(a_bin_pt, b_bin_pt: INTEGER) return INTEGER is
    begin
        return max(a_bin_pt, b_bin_pt);
    end;
    function integer_bits(a_width, a_bin_pt, b_width, b_bin_pt: INTEGER)
        return INTEGER is
    begin
        return  max(a_width - a_bin_pt, b_width - b_bin_pt);
    end;
    function pad_LSB(inp : std_logic_vector; new_width: integer)
        return STD_LOGIC_VECTOR
    is
        constant orig_width : integer := inp'length;
        variable vec : std_logic_vector(orig_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable pos : integer;
        constant pad_pos : integer := new_width - orig_width - 1;
    begin
        vec := inp;
        pos := new_width-1;
        if (new_width >= orig_width) then
            for i in orig_width-1 downto 0 loop
                result(pos) := vec(i);
                pos := pos - 1;
            end loop;
            if pad_pos >= 0 then
                for i in pad_pos downto 0 loop
                    result(i) := '0';
                end loop;
            end if;
        end if;
        return result;
    end;
    function sign_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector
    is
        constant old_width : integer := inp'length;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if new_width >= old_width then
            result(old_width-1 downto 0) := vec;
            if new_width-1 >= old_width then
                for i in new_width-1 downto old_width loop
                    result(i) := vec(old_width-1);
                end loop;
            end if;
        else
            result(new_width-1 downto 0) := vec(new_width-1 downto 0);
        end if;
        return result;
    end;
    function zero_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector
    is
        constant old_width : integer := inp'length;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if new_width >= old_width then
            result(old_width-1 downto 0) := vec;
            if new_width-1 >= old_width then
                for i in new_width-1 downto old_width loop
                    result(i) := '0';
                end loop;
            end if;
        else
            result(new_width-1 downto 0) := vec(new_width-1 downto 0);
        end if;
        return result;
    end;
    function zero_ext(inp : std_logic; new_width : INTEGER)
        return std_logic_vector
    is
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        result(0) := inp;
        for i in new_width-1 downto 1 loop
            result(i) := '0';
        end loop;
        return result;
    end;
    function extend_MSB(inp : std_logic_vector; new_width, arith : INTEGER)
        return std_logic_vector
    is
        constant orig_width : integer := inp'length;
        variable vec : std_logic_vector(orig_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if arith = xlUnsigned then
            result := zero_ext(vec, new_width);
        else
            result := sign_ext(vec, new_width);
        end if;
        return result;
    end;
    function pad_LSB(inp : std_logic_vector; new_width, arith: integer)
        return STD_LOGIC_VECTOR
    is
        constant orig_width : integer := inp'length;
        variable vec : std_logic_vector(orig_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable pos : integer;
    begin
        vec := inp;
        pos := new_width-1;
        if (arith = xlUnsigned) then
            result(pos) := '0';
            pos := pos - 1;
        else
            result(pos) := vec(orig_width-1);
            pos := pos - 1;
        end if;
        if (new_width >= orig_width) then
            for i in orig_width-1 downto 0 loop
                result(pos) := vec(i);
                pos := pos - 1;
            end loop;
            if pos >= 0 then
                for i in pos downto 0 loop
                    result(i) := '0';
                end loop;
            end if;
        end if;
        return result;
    end;
    function align_input(inp : std_logic_vector; old_width, delta, new_arith,
                         new_width: INTEGER)
        return std_logic_vector
    is
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable padded_inp : std_logic_vector((old_width + delta)-1  downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if delta > 0 then
            padded_inp := pad_LSB(vec, old_width+delta);
            result := extend_MSB(padded_inp, new_width, new_arith);
        else
            result := extend_MSB(vec, new_width, new_arith);
        end if;
        return result;
    end;
    function max(L, R: INTEGER) return INTEGER is
    begin
        if L > R then
            return L;
        else
            return R;
        end if;
    end;
    function min(L, R: INTEGER) return INTEGER is
    begin
        if L < R then
            return L;
        else
            return R;
        end if;
    end;
    function "="(left,right: STRING) return boolean is
    begin
        if (left'length /= right'length) then
            return false;
        else
            test : for i in 1 to left'length loop
                if left(i) /= right(i) then
                    return false;
                end if;
            end loop test;
            return true;
        end if;
    end;
    -- synopsys translate_off
    function is_binary_string_invalid (inp : string)
        return boolean
    is
        variable vec : string(1 to inp'length);
        variable result : boolean;
    begin
        vec := inp;
        result := false;
        for i in 1 to vec'length loop
            if ( vec(i) = 'X' ) then
                result := true;
            end if;
        end loop;
        return result;
    end;
    function is_binary_string_undefined (inp : string)
        return boolean
    is
        variable vec : string(1 to inp'length);
        variable result : boolean;
    begin
        vec := inp;
        result := false;
        for i in 1 to vec'length loop
            if ( vec(i) = 'U' ) then
                result := true;
            end if;
        end loop;
        return result;
    end;
    function is_XorU(inp : std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        vec := inp;
        result := false;
        for i in 0 to width-1 loop
            if (vec(i) = 'U') or (vec(i) = 'X') then
                result := true;
            end if;
        end loop;
        return result;
    end;
    function to_real(inp : std_logic_vector; bin_pt : integer; arith : integer)
        return real
    is
        variable  vec : std_logic_vector(inp'length-1 downto 0);
        variable result, shift_val, undefined_real : real;
        variable neg_num : boolean;
    begin
        vec := inp;
        result := 0.0;
        neg_num := false;
        if vec(inp'length-1) = '1' then
            neg_num := true;
        end if;
        for i in 0 to inp'length-1 loop
            if  vec(i) = 'U' or vec(i) = 'X' then
                return undefined_real;
            end if;
            if arith = xlSigned then
                if neg_num then
                    if vec(i) = '0' then
                        result := result + 2.0**i;
                    end if;
                else
                    if vec(i) = '1' then
                        result := result + 2.0**i;
                    end if;
                end if;
            else
                if vec(i) = '1' then
                    result := result + 2.0**i;
                end if;
            end if;
        end loop;
        if arith = xlSigned then
            if neg_num then
                result := result + 1.0;
                result := result * (-1.0);
            end if;
        end if;
        shift_val := 2.0**(-1*bin_pt);
        result := result * shift_val;
        return result;
    end;
    function std_logic_to_real(inp : std_logic; bin_pt : integer; arith : integer)
        return real
    is
        variable result : real := 0.0;
    begin
        if inp = '1' then
            result := 1.0;
        end if;
        if arith = xlSigned then
            assert false
                report "It doesn't make sense to convert a 1 bit number to a signed real.";
        end if;
        return result;
    end;
    -- synopsys translate_on
    function integer_to_std_logic_vector (inp : integer;  width, arith : integer)
        return std_logic_vector
    is
        variable result : std_logic_vector(width-1 downto 0);
        variable unsigned_val : unsigned(width-1 downto 0);
        variable signed_val : signed(width-1 downto 0);
    begin
        if (arith = xlSigned) then
            signed_val := to_signed(inp, width);
            result := signed_to_std_logic_vector(signed_val);
        else
            unsigned_val := to_unsigned(inp, width);
            result := unsigned_to_std_logic_vector(unsigned_val);
        end if;
        return result;
    end;
    function std_logic_vector_to_integer (inp : std_logic_vector;  arith : integer)
        return integer
    is
        constant width : integer := inp'length;
        variable unsigned_val : unsigned(width-1 downto 0);
        variable signed_val : signed(width-1 downto 0);
        variable result : integer;
    begin
        if (arith = xlSigned) then
            signed_val := std_logic_vector_to_signed(inp);
            result := to_integer(signed_val);
        else
            unsigned_val := std_logic_vector_to_unsigned(inp);
            result := to_integer(unsigned_val);
        end if;
        return result;
    end;
    function std_logic_to_integer(constant inp : std_logic := '0')
        return integer
    is
    begin
        if inp = '1' then
            return 1;
        else
            return 0;
        end if;
    end;
    function makeZeroBinStr (width : integer) return STRING is
        variable result : string(1 to width+3);
    begin
        result(1) := '0';
        result(2) := 'b';
        for i in 3 to width+2 loop
            result(i) := '0';
        end loop;
        result(width+3) := '.';
        return result;
    end;
    -- synopsys translate_off
    function real_string_to_std_logic_vector (inp : string;  width, bin_pt, arith : integer)
        return std_logic_vector
    is
        variable result : std_logic_vector(width-1 downto 0);
    begin
        result := (others => '0');
        return result;
    end;
    function real_to_std_logic_vector (inp : real;  width, bin_pt, arith : integer)
        return std_logic_vector
    is
        variable real_val : real;
        variable int_val : integer;
        variable result : std_logic_vector(width-1 downto 0) := (others => '0');
        variable unsigned_val : unsigned(width-1 downto 0) := (others => '0');
        variable signed_val : signed(width-1 downto 0) := (others => '0');
    begin
        real_val := inp;
        int_val := integer(real_val * 2.0**(bin_pt));
        if (arith = xlSigned) then
            signed_val := to_signed(int_val, width);
            result := signed_to_std_logic_vector(signed_val);
        else
            unsigned_val := to_unsigned(int_val, width);
            result := unsigned_to_std_logic_vector(unsigned_val);
        end if;
        return result;
    end;
    -- synopsys translate_on
    function valid_bin_string (inp : string)
        return boolean
    is
        variable vec : string(1 to inp'length);
    begin
        vec := inp;
        if (vec(1) = '0' and vec(2) = 'b') then
            return true;
        else
            return false;
        end if;
    end;
    function hex_string_to_std_logic_vector(inp: string; width : integer)
        return std_logic_vector is
        constant strlen       : integer := inp'LENGTH;
        variable result       : std_logic_vector(width-1 downto 0);
        variable bitval       : std_logic_vector((strlen*4)-1 downto 0);
        variable posn         : integer;
        variable ch           : character;
        variable vec          : string(1 to strlen);
    begin
        vec := inp;
        result := (others => '0');
        posn := (strlen*4)-1;
        for i in 1 to strlen loop
            ch := vec(i);
            case ch is
                when '0' => bitval(posn downto posn-3) := "0000";
                when '1' => bitval(posn downto posn-3) := "0001";
                when '2' => bitval(posn downto posn-3) := "0010";
                when '3' => bitval(posn downto posn-3) := "0011";
                when '4' => bitval(posn downto posn-3) := "0100";
                when '5' => bitval(posn downto posn-3) := "0101";
                when '6' => bitval(posn downto posn-3) := "0110";
                when '7' => bitval(posn downto posn-3) := "0111";
                when '8' => bitval(posn downto posn-3) := "1000";
                when '9' => bitval(posn downto posn-3) := "1001";
                when 'A' | 'a' => bitval(posn downto posn-3) := "1010";
                when 'B' | 'b' => bitval(posn downto posn-3) := "1011";
                when 'C' | 'c' => bitval(posn downto posn-3) := "1100";
                when 'D' | 'd' => bitval(posn downto posn-3) := "1101";
                when 'E' | 'e' => bitval(posn downto posn-3) := "1110";
                when 'F' | 'f' => bitval(posn downto posn-3) := "1111";
                when others => bitval(posn downto posn-3) := "XXXX";
                               -- synopsys translate_off
                               ASSERT false
                                   REPORT "Invalid hex value" SEVERITY ERROR;
                               -- synopsys translate_on
            end case;
            posn := posn - 4;
        end loop;
        if (width <= strlen*4) then
            result :=  bitval(width-1 downto 0);
        else
            result((strlen*4)-1 downto 0) := bitval;
        end if;
        return result;
    end;
    function bin_string_to_std_logic_vector (inp : string)
        return std_logic_vector
    is
        variable pos : integer;
        variable vec : string(1 to inp'length);
        variable result : std_logic_vector(inp'length-1 downto 0);
    begin
        vec := inp;
        pos := inp'length-1;
        result := (others => '0');
        for i in 1 to vec'length loop
            -- synopsys translate_off
            if (pos < 0) and (vec(i) = '0' or vec(i) = '1' or vec(i) = 'X' or vec(i) = 'U')  then
                assert false
                    report "Input string is larger than output std_logic_vector. Truncating output.";
                return result;
            end if;
            -- synopsys translate_on
            if vec(i) = '0' then
                result(pos) := '0';
                pos := pos - 1;
            end if;
            if vec(i) = '1' then
                result(pos) := '1';
                pos := pos - 1;
            end if;
            -- synopsys translate_off
            if (vec(i) = 'X' or vec(i) = 'U') then
                result(pos) := 'U';
                pos := pos - 1;
            end if;
            -- synopsys translate_on
        end loop;
        return result;
    end;
    function bin_string_element_to_std_logic_vector (inp : string;  width, index : integer)
        return std_logic_vector
    is
        constant str_width : integer := width + 4;
        constant inp_len : integer := inp'length;
        constant num_elements : integer := (inp_len + 1)/str_width;
        constant reverse_index : integer := (num_elements-1) - index;
        variable left_pos : integer;
        variable right_pos : integer;
        variable vec : string(1 to inp'length);
        variable result : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        result := (others => '0');
        if (reverse_index = 0) and (reverse_index < num_elements) and (inp_len-3 >= width) then
            left_pos := 1;
            right_pos := width + 3;
            result := bin_string_to_std_logic_vector(vec(left_pos to right_pos));
        end if;
        if (reverse_index > 0) and (reverse_index < num_elements) and (inp_len-3 >= width) then
            left_pos := (reverse_index * str_width) + 1;
            right_pos := left_pos + width + 2;
            result := bin_string_to_std_logic_vector(vec(left_pos to right_pos));
        end if;
        return result;
    end;
   -- synopsys translate_off
    function std_logic_vector_to_bin_string(inp : std_logic_vector)
        return string
    is
        variable vec : std_logic_vector(1 to inp'length);
        variable result : string(vec'range);
    begin
        vec := inp;
        for i in vec'range loop
            result(i) := to_char(vec(i));
        end loop;
        return result;
    end;
    function std_logic_to_bin_string(inp : std_logic)
        return string
    is
        variable result : string(1 to 3);
    begin
        result(1) := '0';
        result(2) := 'b';
        result(3) := to_char(inp);
        return result;
    end;
    function std_logic_vector_to_bin_string_w_point(inp : std_logic_vector; bin_pt : integer)
        return string
    is
        variable width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable str_pos : integer;
        variable result : string(1 to width+3);
    begin
        vec := inp;
        str_pos := 1;
        result(str_pos) := '0';
        str_pos := 2;
        result(str_pos) := 'b';
        str_pos := 3;
        for i in width-1 downto 0  loop
            if (((width+3) - bin_pt) = str_pos) then
                result(str_pos) := '.';
                str_pos := str_pos + 1;
            end if;
            result(str_pos) := to_char(vec(i));
            str_pos := str_pos + 1;
        end loop;
        if (bin_pt = 0) then
            result(str_pos) := '.';
        end if;
        return result;
    end;
    function real_to_bin_string(inp : real;  width, bin_pt, arith : integer)
        return string
    is
        variable result : string(1 to width);
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := real_to_std_logic_vector(inp, width, bin_pt, arith);
        result := std_logic_vector_to_bin_string(vec);
        return result;
    end;
    function real_to_string (inp : real) return string
    is
        variable result : string(1 to display_precision) := (others => ' ');
    begin
        result(real'image(inp)'range) := real'image(inp);
        return result;
    end;
    -- synopsys translate_on
end conv_pkg;

-------------------------------------------------------------------
-- System Generator version 13.2 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
library warp_per_block_calc_lib;
use warp_per_block_calc_lib.conv_pkg.all;
entity srl17e is
    generic (width : integer:=16;
             latency : integer :=8);
    port (clk   : in std_logic;
          ce    : in std_logic;
          d     : in std_logic_vector(width-1 downto 0);
          q     : out std_logic_vector(width-1 downto 0));
end srl17e;
architecture structural of srl17e is
    component SRL16E
        port (D   : in STD_ULOGIC;
              CE  : in STD_ULOGIC;
              CLK : in STD_ULOGIC;
              A0  : in STD_ULOGIC;
              A1  : in STD_ULOGIC;
              A2  : in STD_ULOGIC;
              A3  : in STD_ULOGIC;
              Q   : out STD_ULOGIC);
    end component;
    attribute syn_black_box of SRL16E : component is true;
    attribute fpga_dont_touch of SRL16E : component is "true";
    component FDE
        port(
            Q  :        out   STD_ULOGIC;
            D  :        in    STD_ULOGIC;
            C  :        in    STD_ULOGIC;
            CE :        in    STD_ULOGIC);
    end component;
    attribute syn_black_box of FDE : component is true;
    attribute fpga_dont_touch of FDE : component is "true";
    constant a : std_logic_vector(4 downto 0) :=
        integer_to_std_logic_vector(latency-2,5,xlSigned);
    signal d_delayed : std_logic_vector(width-1 downto 0);
    signal srl16_out : std_logic_vector(width-1 downto 0);
begin
    d_delayed <= d after 200 ps;
    reg_array : for i in 0 to width-1 generate
        srl16_used: if latency > 1 generate
            u1 : srl16e port map(clk => clk,
                                 d => d_delayed(i),
                                 q => srl16_out(i),
                                 ce => ce,
                                 a0 => a(0),
                                 a1 => a(1),
                                 a2 => a(2),
                                 a3 => a(3));
        end generate;
        srl16_not_used: if latency <= 1 generate
            srl16_out(i) <= d_delayed(i);
        end generate;
        fde_used: if latency /= 0  generate
            u2 : fde port map(c => clk,
                              d => srl16_out(i),
                              q => q(i),
                              ce => ce);
        end generate;
        fde_not_used: if latency = 0  generate
            q(i) <= srl16_out(i);
        end generate;
    end generate;
 end structural;
library IEEE;
use IEEE.std_logic_1164.all;
library warp_per_block_calc_lib;
use warp_per_block_calc_lib.conv_pkg.all;
entity synth_reg is
    generic (width           : integer := 8;
             latency         : integer := 1);
    port (i       : in std_logic_vector(width-1 downto 0);
          ce      : in std_logic;
          clr     : in std_logic;
          clk     : in std_logic;
          o       : out std_logic_vector(width-1 downto 0));
end synth_reg;
architecture structural of synth_reg is
    component srl17e
        generic (width : integer:=16;
                 latency : integer :=8);
        port (clk : in std_logic;
              ce  : in std_logic;
              d   : in std_logic_vector(width-1 downto 0);
              q   : out std_logic_vector(width-1 downto 0));
    end component;
    function calc_num_srl17es (latency : integer)
        return integer
    is
        variable remaining_latency : integer;
        variable result : integer;
    begin
        result := latency / 17;
        remaining_latency := latency - (result * 17);
        if (remaining_latency /= 0) then
            result := result + 1;
        end if;
        return result;
    end;
    constant complete_num_srl17es : integer := latency / 17;
    constant num_srl17es : integer := calc_num_srl17es(latency);
    constant remaining_latency : integer := latency - (complete_num_srl17es * 17);
    type register_array is array (num_srl17es downto 0) of
        std_logic_vector(width-1 downto 0);
    signal z : register_array;
begin
    z(0) <= i;
    complete_ones : if complete_num_srl17es > 0 generate
        srl17e_array: for i in 0 to complete_num_srl17es-1 generate
            delay_comp : srl17e
                generic map (width => width,
                             latency => 17)
                port map (clk => clk,
                          ce  => ce,
                          d       => z(i),
                          q       => z(i+1));
        end generate;
    end generate;
    partial_one : if remaining_latency > 0 generate
        last_srl17e : srl17e
            generic map (width => width,
                         latency => remaining_latency)
            port map (clk => clk,
                      ce  => ce,
                      d   => z(num_srl17es-1),
                      q   => z(num_srl17es));
    end generate;
    o <= z(num_srl17es);
end structural;
library IEEE;
use IEEE.std_logic_1164.all;
library warp_per_block_calc_lib;
use warp_per_block_calc_lib.conv_pkg.all;
entity synth_reg_reg is
    generic (width           : integer := 8;
             latency         : integer := 1);
    port (i       : in std_logic_vector(width-1 downto 0);
          ce      : in std_logic;
          clr     : in std_logic;
          clk     : in std_logic;
          o       : out std_logic_vector(width-1 downto 0));
end synth_reg_reg;
architecture behav of synth_reg_reg is
  type reg_array_type is array (latency-1 downto 0) of std_logic_vector(width -1 downto 0);
  signal reg_bank : reg_array_type := (others => (others => '0'));
  signal reg_bank_in : reg_array_type := (others => (others => '0'));
  attribute syn_allow_retiming : boolean;
  attribute syn_srlstyle : string;
  attribute syn_allow_retiming of reg_bank : signal is true;
  attribute syn_allow_retiming of reg_bank_in : signal is true;
  attribute syn_srlstyle of reg_bank : signal is "registers";
  attribute syn_srlstyle of reg_bank_in : signal is "registers";
begin
  latency_eq_0: if latency = 0 generate
    o <= i;
  end generate latency_eq_0;
  latency_gt_0: if latency >= 1 generate
    o <= reg_bank(latency-1);
    reg_bank_in(0) <= i;
    loop_gen: for idx in latency-2 downto 0 generate
      reg_bank_in(idx+1) <= reg_bank(idx);
    end generate loop_gen;
    sync_loop: for sync_idx in latency-1 downto 0 generate
      sync_proc: process (clk)
      begin
        if clk'event and clk = '1' then
          if ce = '1'  then
            reg_bank(sync_idx) <= reg_bank_in(sync_idx);
          end if;
        end if;
      end process sync_proc;
    end generate sync_loop;
  end generate latency_gt_0;
end behav;

-------------------------------------------------------------------
-- System Generator version 13.2 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
library warp_per_block_calc_lib;
use warp_per_block_calc_lib.conv_pkg.all;
entity single_reg_w_init is
  generic (
    width: integer := 8;
    init_index: integer := 0;
    init_value: bit_vector := b"0000"
  );
  port (
    i: in std_logic_vector(width - 1 downto 0);
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    o: out std_logic_vector(width - 1 downto 0)
  );
end single_reg_w_init;
architecture structural of single_reg_w_init is
  function build_init_const(width: integer;
                            init_index: integer;
                            init_value: bit_vector)
    return std_logic_vector
  is
    variable result: std_logic_vector(width - 1 downto 0);
  begin
    if init_index = 0 then
      result := (others => '0');
    elsif init_index = 1 then
      result := (others => '0');
      result(0) := '1';
    else
      result := to_stdlogicvector(init_value);
    end if;
    return result;
  end;
  component fdre
    port (
      q: out std_ulogic;
      d: in  std_ulogic;
      c: in  std_ulogic;
      ce: in  std_ulogic;
      r: in  std_ulogic
    );
  end component;
  attribute syn_black_box of fdre: component is true;
  attribute fpga_dont_touch of fdre: component is "true";
  component fdse
    port (
      q: out std_ulogic;
      d: in  std_ulogic;
      c: in  std_ulogic;
      ce: in  std_ulogic;
      s: in  std_ulogic
    );
  end component;
  attribute syn_black_box of fdse: component is true;
  attribute fpga_dont_touch of fdse: component is "true";
  constant init_const: std_logic_vector(width - 1 downto 0)
    := build_init_const(width, init_index, init_value);
begin
  fd_prim_array: for index in 0 to width - 1 generate
    bit_is_0: if (init_const(index) = '0') generate
      fdre_comp: fdre
        port map (
          c => clk,
          d => i(index),
          q => o(index),
          ce => ce,
          r => clr
        );
    end generate;
    bit_is_1: if (init_const(index) = '1') generate
      fdse_comp: fdse
        port map (
          c => clk,
          d => i(index),
          q => o(index),
          ce => ce,
          s => clr
        );
    end generate;
  end generate;
end architecture structural;
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
library warp_per_block_calc_lib;
use warp_per_block_calc_lib.conv_pkg.all;
entity synth_reg_w_init is
  generic (
    width: integer := 8;
    init_index: integer := 0;
    init_value: bit_vector := b"0000";
    latency: integer := 1
  );
  port (
    i: in std_logic_vector(width - 1 downto 0);
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    o: out std_logic_vector(width - 1 downto 0)
  );
end synth_reg_w_init;
architecture structural of synth_reg_w_init is
  component single_reg_w_init
    generic (
      width: integer := 8;
      init_index: integer := 0;
      init_value: bit_vector := b"0000"
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  signal dly_i: std_logic_vector((latency + 1) * width - 1 downto 0);
  signal dly_clr: std_logic;
begin
  latency_eq_0: if (latency = 0) generate
    o <= i;
  end generate;
  latency_gt_0: if (latency >= 1) generate
    dly_i((latency + 1) * width - 1 downto latency * width) <= i
      after 200 ps;
    dly_clr <= clr after 200 ps;
    fd_array: for index in latency downto 1 generate
       reg_comp: single_reg_w_init
          generic map (
            width => width,
            init_index => init_index,
            init_value => init_value
          )
          port map (
            clk => clk,
            i => dly_i((index + 1) * width - 1 downto index * width),
            o => dly_i(index * width - 1 downto (index - 1) * width),
            ce => ce,
            clr => dly_clr
          );
    end generate;
    o <= dly_i(width - 1 downto 0);
  end generate;
end structural;

-------------------------------------------------------------------
-- System Generator version 13.2 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
library warp_per_block_calc_lib;
use warp_per_block_calc_lib.conv_pkg.all;
entity xladdsub is
  generic (
    core_name0: string := "";
    a_width: integer := 16;
    a_bin_pt: integer := 4;
    a_arith: integer := xlUnsigned;
    c_in_width: integer := 16;
    c_in_bin_pt: integer := 4;
    c_in_arith: integer := xlUnsigned;
    c_out_width: integer := 16;
    c_out_bin_pt: integer := 4;
    c_out_arith: integer := xlUnsigned;
    b_width: integer := 8;
    b_bin_pt: integer := 2;
    b_arith: integer := xlUnsigned;
    s_width: integer := 17;
    s_bin_pt: integer := 4;
    s_arith: integer := xlUnsigned;
    rst_width: integer := 1;
    rst_bin_pt: integer := 0;
    rst_arith: integer := xlUnsigned;
    en_width: integer := 1;
    en_bin_pt: integer := 0;
    en_arith: integer := xlUnsigned;
    full_s_width: integer := 17;
    full_s_arith: integer := xlUnsigned;
    mode: integer := xlAddMode;
    extra_registers: integer := 0;
    latency: integer := 0;
    quantization: integer := xlTruncate;
    overflow: integer := xlWrap;
    c_latency: integer := 0;
    c_output_width: integer := 17;
    c_has_c_in : integer := 0;
    c_has_c_out : integer := 0
  );
  port (
    a: in std_logic_vector(a_width - 1 downto 0);
    b: in std_logic_vector(b_width - 1 downto 0);
    c_in : in std_logic_vector (0 downto 0) := "0";
    ce: in std_logic;
    clr: in std_logic := '0';
    clk: in std_logic;
    rst: in std_logic_vector(rst_width - 1 downto 0) := "0";
    en: in std_logic_vector(en_width - 1 downto 0) := "1";
    c_out : out std_logic_vector (0 downto 0);
    s: out std_logic_vector(s_width - 1 downto 0)
  );
end xladdsub;
architecture behavior of xladdsub is
  component synth_reg
    generic (
      width: integer := 16;
      latency: integer := 5
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  function format_input(inp: std_logic_vector; old_width, delta, new_arith,
                        new_width: integer)
    return std_logic_vector
  is
    variable vec: std_logic_vector(old_width-1 downto 0);
    variable padded_inp: std_logic_vector((old_width + delta)-1  downto 0);
    variable result: std_logic_vector(new_width-1 downto 0);
  begin
    vec := inp;
    if (delta > 0) then
      padded_inp := pad_LSB(vec, old_width+delta);
      result := extend_MSB(padded_inp, new_width, new_arith);
    else
      result := extend_MSB(vec, new_width, new_arith);
    end if;
    return result;
  end;
  constant full_s_bin_pt: integer := fractional_bits(a_bin_pt, b_bin_pt);
  constant full_a_width: integer := full_s_width;
  constant full_b_width: integer := full_s_width;
  signal full_a: std_logic_vector(full_a_width - 1 downto 0);
  signal full_b: std_logic_vector(full_b_width - 1 downto 0);
  signal core_s: std_logic_vector(full_s_width - 1 downto 0);
  signal conv_s: std_logic_vector(s_width - 1 downto 0);
  signal temp_cout : std_logic;
  signal internal_clr: std_logic;
  signal internal_ce: std_logic;
  signal extra_reg_ce: std_logic;
  signal override: std_logic;
  signal logic1: std_logic_vector(0 downto 0);
  component addsb_11_0_84fc5d4200208b4e
    port (
          a: in std_logic_vector(7 - 1 downto 0);
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(7 - 1 downto 0)
    );
  end component;
  attribute syn_black_box of addsb_11_0_84fc5d4200208b4e:
    component is true;
  attribute fpga_dont_touch of addsb_11_0_84fc5d4200208b4e:
    component is "true";
  attribute box_type of addsb_11_0_84fc5d4200208b4e:
    component  is "black_box";
begin
  internal_clr <= (clr or (rst(0))) and ce;
  internal_ce <= ce and en(0);
  logic1(0) <= '1';
  addsub_process: process (a, b, core_s)
  begin
    full_a <= format_input (a, a_width, b_bin_pt - a_bin_pt, a_arith,
                            full_a_width);
    full_b <= format_input (b, b_width, a_bin_pt - b_bin_pt, b_arith,
                            full_b_width);
    conv_s <= convert_type (core_s, full_s_width, full_s_bin_pt, full_s_arith,
                            s_width, s_bin_pt, s_arith, quantization, overflow);
  end process addsub_process;

  comp0: if ((core_name0 = "addsb_11_0_84fc5d4200208b4e")) generate
    core_instance0: addsb_11_0_84fc5d4200208b4e
      port map (
         a => full_a,
         s => core_s,
         b => full_b
      );
  end generate;
  latency_test: if (extra_registers > 0) generate
      override_test: if (c_latency > 1) generate
       override_pipe: synth_reg
          generic map (
            width => 1,
            latency => c_latency
          )
          port map (
            i => logic1,
            ce => internal_ce,
            clr => internal_clr,
            clk => clk,
            o(0) => override);
       extra_reg_ce <= ce and en(0) and override;
      end generate override_test;
      no_override: if ((c_latency = 0) or (c_latency = 1)) generate
       extra_reg_ce <= ce and en(0);
      end generate no_override;
      extra_reg: synth_reg
        generic map (
          width => s_width,
          latency => extra_registers
        )
        port map (
          i => conv_s,
          ce => extra_reg_ce,
          clr => internal_clr,
          clk => clk,
          o => s
        );
      cout_test: if (c_has_c_out = 1) generate
      c_out_extra_reg: synth_reg
        generic map (
          width => 1,
          latency => extra_registers
        )
        port map (
          i(0) => temp_cout,
          ce => extra_reg_ce,
          clr => internal_clr,
          clk => clk,
          o => c_out
        );
      end generate cout_test;
  end generate;
  latency_s: if ((latency = 0) or (extra_registers = 0)) generate
    s <= conv_s;
  end generate latency_s;
  latency0: if (((latency = 0) or (extra_registers = 0)) and
                 (c_has_c_out = 1)) generate
    c_out(0) <= temp_cout;
  end generate latency0;
  tie_dangling_cout: if (c_has_c_out = 0) generate
    c_out <= "0";
  end generate tie_dangling_cout;
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library warp_per_block_calc_lib;
use warp_per_block_calc_lib.conv_pkg.all;

entity constant_963ed6358a is
  port (
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_963ed6358a;


architecture behavior of constant_963ed6358a is
begin
  op <= "0";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library warp_per_block_calc_lib;
use warp_per_block_calc_lib.conv_pkg.all;

entity constant_8567b21c7f is
  port (
    op : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_8567b21c7f;


architecture behavior of constant_8567b21c7f is
begin
  op <= "00100000";
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library warp_per_block_calc_lib;
use warp_per_block_calc_lib.conv_pkg.all;

entity constant_a267c870be is
  port (
    op : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_a267c870be;


architecture behavior of constant_a267c870be is
begin
  op <= "000001";
end behavior;


-------------------------------------------------------------------
-- System Generator version 13.2 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
library warp_per_block_calc_lib;
use warp_per_block_calc_lib.conv_pkg.all;
entity convert_func_call is
    generic (
        din_width    : integer := 16;
        din_bin_pt   : integer := 4;
        din_arith    : integer := xlUnsigned;
        dout_width   : integer := 8;
        dout_bin_pt  : integer := 2;
        dout_arith   : integer := xlUnsigned;
        quantization : integer := xlTruncate;
        overflow     : integer := xlWrap);
    port (
        din : in std_logic_vector (din_width-1 downto 0);
        result : out std_logic_vector (dout_width-1 downto 0));
end convert_func_call;
architecture behavior of convert_func_call is
begin
    result <= convert_type(din, din_width, din_bin_pt, din_arith,
                           dout_width, dout_bin_pt, dout_arith,
                           quantization, overflow);
end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library warp_per_block_calc_lib;
use warp_per_block_calc_lib.conv_pkg.all;
entity xlconvert is
    generic (
        din_width    : integer := 16;
        din_bin_pt   : integer := 4;
        din_arith    : integer := xlUnsigned;
        dout_width   : integer := 8;
        dout_bin_pt  : integer := 2;
        dout_arith   : integer := xlUnsigned;
        en_width     : integer := 1;
        en_bin_pt    : integer := 0;
        en_arith     : integer := xlUnsigned;
        bool_conversion : integer :=0;
        latency      : integer := 0;
        quantization : integer := xlTruncate;
        overflow     : integer := xlWrap);
    port (
        din : in std_logic_vector (din_width-1 downto 0);
        en  : in std_logic_vector (en_width-1 downto 0);
        ce  : in std_logic;
        clr : in std_logic;
        clk : in std_logic;
        dout : out std_logic_vector (dout_width-1 downto 0));
end xlconvert;
architecture behavior of xlconvert is
    component synth_reg
        generic (width       : integer;
                 latency     : integer);
        port (i       : in std_logic_vector(width-1 downto 0);
              ce      : in std_logic;
              clr     : in std_logic;
              clk     : in std_logic;
              o       : out std_logic_vector(width-1 downto 0));
    end component;
    component convert_func_call
        generic (
            din_width    : integer := 16;
            din_bin_pt   : integer := 4;
            din_arith    : integer := xlUnsigned;
            dout_width   : integer := 8;
            dout_bin_pt  : integer := 2;
            dout_arith   : integer := xlUnsigned;
            quantization : integer := xlTruncate;
            overflow     : integer := xlWrap);
        port (
            din : in std_logic_vector (din_width-1 downto 0);
            result : out std_logic_vector (dout_width-1 downto 0));
    end component;
    -- synopsys translate_off
    -- synopsys translate_on
    signal result : std_logic_vector(dout_width-1 downto 0);
    signal internal_ce : std_logic;
begin
    -- synopsys translate_off
    -- synopsys translate_on
    internal_ce <= ce and en(0);

    bool_conversion_generate : if (bool_conversion = 1)
    generate
      result <= din;
    end generate;
    std_conversion_generate : if (bool_conversion = 0)
    generate
      convert : convert_func_call
        generic map (
          din_width   => din_width,
          din_bin_pt  => din_bin_pt,
          din_arith   => din_arith,
          dout_width  => dout_width,
          dout_bin_pt => dout_bin_pt,
          dout_arith  => dout_arith,
          quantization => quantization,
          overflow     => overflow)
        port map (
          din => din,
          result => result);
    end generate;
    latency_test : if (latency > 0) generate
        reg : synth_reg
            generic map (
              width => dout_width,
              latency => latency
            )
            port map (
              i => result,
              ce => internal_ce,
              clr => clr,
              clk => clk,
              o => dout
            );
    end generate;
    latency0 : if (latency = 0)
    generate
        dout <= result;
    end generate latency0;
end  behavior;

-------------------------------------------------------------------
-- System Generator version 13.2 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
library warp_per_block_calc_lib;
use warp_per_block_calc_lib.conv_pkg.all;
entity xlcounter_free is
  generic (
    core_name0: string := "";
    op_width: integer := 5;
    op_arith: integer := xlSigned
  );
  port (
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    op: out std_logic_vector(op_width - 1 downto 0);
    up: in std_logic_vector(0 downto 0) := (others => '0');
    load: in std_logic_vector(0 downto 0) := (others => '0');
    din: in std_logic_vector(op_width - 1 downto 0) := (others => '0');
    en: in std_logic_vector(0 downto 0);
    rst: in std_logic_vector(0 downto 0)
  );
end xlcounter_free ;
architecture behavior of xlcounter_free is
  component cntr_11_0_e7514e290b172ea1
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;
  attribute syn_black_box of cntr_11_0_e7514e290b172ea1:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_e7514e290b172ea1:
    component is "true";
  attribute box_type of cntr_11_0_e7514e290b172ea1:
    component  is "black_box";
-- synopsys translate_off
  constant zeroVec: std_logic_vector(op_width - 1 downto 0) := (others => '0');
  constant oneVec: std_logic_vector(op_width - 1 downto 0) := (others => '1');
  constant zeroStr: string(1 to op_width) :=
    std_logic_vector_to_bin_string(zeroVec);
  constant oneStr: string(1 to op_width) :=
    std_logic_vector_to_bin_string(oneVec);
-- synopsys translate_on
  signal core_sinit: std_logic;
  signal core_ce: std_logic;
  signal op_net: std_logic_vector(op_width - 1 downto 0);
begin
  core_ce <= ce and en(0);
  core_sinit <= (clr or rst(0)) and ce;
  op <= op_net;
  comp0: if ((core_name0 = "cntr_11_0_e7514e290b172ea1")) generate
    core_instance0: cntr_11_0_e7514e290b172ea1
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
end behavior;

-------------------------------------------------------------------
-- System Generator version 13.2 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
library warp_per_block_calc_lib;
use warp_per_block_calc_lib.conv_pkg.all;
entity xldelay is
   generic(width        : integer := -1;
           latency      : integer := -1;
           reg_retiming : integer := 0);
   port(d       : in std_logic_vector (width-1 downto 0);
        ce      : in std_logic;
        clk     : in std_logic;
        en      : in std_logic;
        q       : out std_logic_vector (width-1 downto 0));
end xldelay;
architecture behavior of xldelay is
   component synth_reg
      generic (width       : integer;
               latency     : integer);
      port (i       : in std_logic_vector(width-1 downto 0);
            ce      : in std_logic;
            clr     : in std_logic;
            clk     : in std_logic;
            o       : out std_logic_vector(width-1 downto 0));
   end component;
   component synth_reg_reg
      generic (width       : integer;
               latency     : integer);
      port (i       : in std_logic_vector(width-1 downto 0);
            ce      : in std_logic;
            clr     : in std_logic;
            clk     : in std_logic;
            o       : out std_logic_vector(width-1 downto 0));
   end component;
   signal internal_ce  : std_logic;
begin
   internal_ce  <= ce and en;
   srl_delay: if (reg_retiming = 0) or (latency < 1) generate
     synth_reg_srl_inst : synth_reg
       generic map (
         width   => width,
         latency => latency)
       port map (
         i   => d,
         ce  => internal_ce,
         clr => '0',
         clk => clk,
         o   => q);
   end generate srl_delay;
   reg_delay: if (reg_retiming = 1) and (latency >= 1) generate
     synth_reg_reg_inst : synth_reg_reg
       generic map (
         width   => width,
         latency => latency)
       port map (
         i   => d,
         ce  => internal_ce,
         clr => '0',
         clk => clk,
         o   => q);
   end generate reg_delay;
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library warp_per_block_calc_lib;
use warp_per_block_calc_lib.conv_pkg.all;

entity xldivider_generator_28bcfda473f2ef787fc4fee0cf6012ce is 
  port(
    ce:in std_logic;
    clk:in std_logic;
    dividend:in std_logic_vector(11 downto 0);
    divisor:in std_logic_vector(5 downto 0);
    fractional:out std_logic_vector(15 downto 0);
    quotient:out std_logic_vector(11 downto 0);
    rfd:out std_logic
  );
end xldivider_generator_28bcfda473f2ef787fc4fee0cf6012ce;


architecture behavior of xldivider_generator_28bcfda473f2ef787fc4fee0cf6012ce  is
  component dv_gn_v3_0_c648497ecac7f882
    port(
      ce:in std_logic;
      clk:in std_logic;
      dividend:in std_logic_vector(11 downto 0);
      divisor:in std_logic_vector(5 downto 0);
      fractional:out std_logic_vector(15 downto 0);
      quotient:out std_logic_vector(11 downto 0);
      rfd:out std_logic
    );
end component;
begin
  dv_gn_v3_0_c648497ecac7f882_instance : dv_gn_v3_0_c648497ecac7f882
    port map(
      ce=>ce,
      clk=>clk,
      dividend=>dividend,
      divisor=>divisor,
      fractional=>fractional,
      quotient=>quotient,
      rfd=>rfd
    );
end  behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library warp_per_block_calc_lib;
use warp_per_block_calc_lib.conv_pkg.all;

entity logical_aacf6e1b0e is
  port (
    d0 : in std_logic_vector((1 - 1) downto 0);
    d1 : in std_logic_vector((1 - 1) downto 0);
    y : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_aacf6e1b0e;


architecture behavior of logical_aacf6e1b0e is
  signal d0_1_24: std_logic;
  signal d1_1_27: std_logic;
  signal fully_2_1_bit: std_logic;
begin
  d0_1_24 <= d0(0);
  d1_1_27 <= d1(0);
  fully_2_1_bit <= d0_1_24 or d1_1_27;
  y <= std_logic_to_vector(fully_2_1_bit);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library warp_per_block_calc_lib;
use warp_per_block_calc_lib.conv_pkg.all;

entity mux_ac2c510b5b is
  port (
    sel : in std_logic_vector((1 - 1) downto 0);
    d0 : in std_logic_vector((6 - 1) downto 0);
    d1 : in std_logic_vector((6 - 1) downto 0);
    y : out std_logic_vector((6 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end mux_ac2c510b5b;


architecture behavior of mux_ac2c510b5b is
  signal sel_1_20: std_logic;
  signal d0_1_24: std_logic_vector((6 - 1) downto 0);
  signal d1_1_27: std_logic_vector((6 - 1) downto 0);
  signal sel_internal_2_1_convert: std_logic_vector((1 - 1) downto 0);
  signal unregy_join_6_1: std_logic_vector((6 - 1) downto 0);
begin
  sel_1_20 <= sel(0);
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  sel_internal_2_1_convert <= cast(std_logic_to_vector(sel_1_20), 0, 1, 0, xlUnsigned);
  proc_switch_6_1: process (d0_1_24, d1_1_27, sel_internal_2_1_convert)
  is
  begin
    case sel_internal_2_1_convert is 
      when "0" =>
        unregy_join_6_1 <= d0_1_24;
      when others =>
        unregy_join_6_1 <= d1_1_27;
    end case;
  end process proc_switch_6_1;
  y <= unregy_join_6_1;
end behavior;


-------------------------------------------------------------------
-- System Generator version 13.2 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
library warp_per_block_calc_lib;
use warp_per_block_calc_lib.conv_pkg.all;
entity xlregister is
   generic (d_width          : integer := 5;
            init_value       : bit_vector := b"00");
   port (d   : in std_logic_vector (d_width-1 downto 0);
         rst : in std_logic_vector(0 downto 0) := "0";
         en  : in std_logic_vector(0 downto 0) := "1";
         ce  : in std_logic;
         clk : in std_logic;
         q   : out std_logic_vector (d_width-1 downto 0));
end xlregister;
architecture behavior of xlregister is
   component synth_reg_w_init
      generic (width      : integer;
               init_index : integer;
               init_value : bit_vector;
               latency    : integer);
      port (i   : in std_logic_vector(width-1 downto 0);
            ce  : in std_logic;
            clr : in std_logic;
            clk : in std_logic;
            o   : out std_logic_vector(width-1 downto 0));
   end component;
   -- synopsys translate_off
   signal real_d, real_q           : real;
   -- synopsys translate_on
   signal internal_clr             : std_logic;
   signal internal_ce              : std_logic;
begin
   internal_clr <= rst(0) and ce;
   internal_ce  <= en(0) and ce;
   synth_reg_inst : synth_reg_w_init
      generic map (width      => d_width,
                   init_index => 2,
                   init_value => init_value,
                   latency    => 1)
      port map (i   => d,
                ce  => internal_ce,
                clr => internal_clr,
                clk => clk,
                o   => q);
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library warp_per_block_calc_lib;
use warp_per_block_calc_lib.conv_pkg.all;

entity relational_54048c8b02 is
  port (
    a : in std_logic_vector((8 - 1) downto 0);
    b : in std_logic_vector((8 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_54048c8b02;


architecture behavior of relational_54048c8b02 is
  signal a_1_31: unsigned((8 - 1) downto 0);
  signal b_1_34: unsigned((8 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library warp_per_block_calc_lib;
use warp_per_block_calc_lib.conv_pkg.all;

entity relational_4eca908438 is
  port (
    a : in std_logic_vector((16 - 1) downto 0);
    b : in std_logic_vector((1 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_4eca908438;


architecture behavior of relational_4eca908438 is
  signal a_1_31: unsigned((16 - 1) downto 0);
  signal b_1_34: unsigned((1 - 1) downto 0);
  signal cast_14_12: unsigned((17 - 1) downto 0);
  signal cast_14_17: unsigned((17 - 1) downto 0);
  signal result_14_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  cast_14_12 <= u2u_cast(a_1_31, 16, 17, 16);
  cast_14_17 <= u2u_cast(b_1_34, 0, 17, 16);
  result_14_3_rel <= cast_14_12 /= cast_14_17;
  op <= boolean_to_vector(result_14_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
library warp_per_block_calc_lib;
use warp_per_block_calc_lib.conv_pkg.all;

-- Generated from Simulink block "warps_per_block_calc"

entity warps_per_block_calc is
  port (
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    en: in std_logic; 
    threads_per_block_in: in std_logic_vector(11 downto 0); 
    warp_size_in: in std_logic_vector(5 downto 0); 
    data_valid_out: out std_logic; 
    warps_per_block_out: out std_logic_vector(5 downto 0)
  );
end warps_per_block_calc;

architecture structural of warps_per_block_calc is
  attribute core_generation_info: string;
  attribute core_generation_info of structural : architecture is "warps_per_block_calc,sysgen_core,{clock_period=10.00000000,clocking=Clock_Enables,compilation=NGC_Netlist,sample_periods=1.00000000000,testbench=1,total_blocks=33,xilinx_adder_subtracter_block=1,xilinx_arithmetic_relational_operator_block=2,xilinx_bus_multiplexer_block=1,xilinx_constant_block_block=3,xilinx_counter_block=1,xilinx_delay_block=1,xilinx_divider_generator_3_0_block=1,xilinx_gateway_in_block=3,xilinx_gateway_out_block=2,xilinx_logical_block_block=1,xilinx_register_block=5,xilinx_resource_estimator_block=1,xilinx_system_generator_block=1,xilinx_type_converter_block=2,}";

  signal addsub_s_net: std_logic_vector(5 downto 0);
  signal ce_1_sg_x0: std_logic;
  signal clk_1_sg_x0: std_logic;
  signal constant1_op_net: std_logic;
  signal constant2_op_net: std_logic_vector(7 downto 0);
  signal constant4_op_net: std_logic_vector(5 downto 0);
  signal convert1_dout_net: std_logic;
  signal convert_dout_net: std_logic_vector(5 downto 0);
  signal counter3_op_net: std_logic_vector(7 downto 0);
  signal data_valid_out_net: std_logic;
  signal delay_q_net: std_logic;
  signal divider_generator_3_0_fractional_net: std_logic_vector(15 downto 0);
  signal divider_generator_3_0_quotient_net: std_logic_vector(11 downto 0);
  signal en_net: std_logic;
  signal logical_y_net: std_logic;
  signal mux_y_net: std_logic_vector(5 downto 0);
  signal register1_q_net: std_logic_vector(11 downto 0);
  signal register3_q_net: std_logic_vector(5 downto 0);
  signal register7_q_net: std_logic;
  signal relational1_op_net: std_logic;
  signal relational_op_net: std_logic;
  signal threads_per_block_in_net: std_logic_vector(11 downto 0);
  signal warp_size_in_net: std_logic_vector(5 downto 0);
  signal warps_per_block_out_net: std_logic_vector(5 downto 0);

begin
  ce_1_sg_x0 <= ce_1;
  clk_1_sg_x0 <= clk_1;
  en_net <= en;
  threads_per_block_in_net <= threads_per_block_in;
  warp_size_in_net <= warp_size_in;
  data_valid_out <= data_valid_out_net;
  warps_per_block_out <= warps_per_block_out_net;

  addsub: entity warp_per_block_calc_lib.xladdsub
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 6,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 6,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 7,
      core_name0 => "addsb_11_0_84fc5d4200208b4e",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 7,
      latency => 0,
      overflow => 1,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 6
    )
    port map (
      a => convert_dout_net,
      b => constant4_op_net,
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      en => "1",
      s => addsub_s_net
    );

  constant1: entity warp_per_block_calc_lib.constant_963ed6358a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => constant1_op_net
    );

  constant2: entity warp_per_block_calc_lib.constant_8567b21c7f
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant2_op_net
    );

  constant4: entity warp_per_block_calc_lib.constant_a267c870be
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant4_op_net
    );

  convert: entity warp_per_block_calc_lib.xlconvert
    generic map (
      bool_conversion => 0,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 12,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 6,
      latency => 0,
      overflow => xlSaturate,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      din => divider_generator_3_0_quotient_net,
      en => "1",
      dout => convert_dout_net
    );

  convert1: entity warp_per_block_calc_lib.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      din(0) => en_net,
      en => "1",
      dout(0) => convert1_dout_net
    );

  counter3: entity warp_per_block_calc_lib.xlcounter_free
    generic map (
      core_name0 => "cntr_11_0_e7514e290b172ea1",
      op_arith => xlUnsigned,
      op_width => 8
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      en(0) => register7_q_net,
      rst(0) => delay_q_net,
      op => counter3_op_net
    );

  delay: entity warp_per_block_calc_lib.xldelay
    generic map (
      latency => 1,
      reg_retiming => 0,
      width => 1
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d(0) => relational_op_net,
      en => '1',
      q(0) => delay_q_net
    );

  divider_generator_3_0: entity warp_per_block_calc_lib.xldivider_generator_28bcfda473f2ef787fc4fee0cf6012ce
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      dividend => register1_q_net,
      divisor => register3_q_net,
      fractional => divider_generator_3_0_fractional_net,
      quotient => divider_generator_3_0_quotient_net
    );

  logical: entity warp_per_block_calc_lib.logical_aacf6e1b0e
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0(0) => relational_op_net,
      d1(0) => convert1_dout_net,
      y(0) => logical_y_net
    );

  mux: entity warp_per_block_calc_lib.mux_ac2c510b5b
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => convert_dout_net,
      d1 => addsub_s_net,
      sel(0) => relational1_op_net,
      y => mux_y_net
    );

  register1: entity warp_per_block_calc_lib.xlregister
    generic map (
      d_width => 12,
      init_value => b"000000000000"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d => threads_per_block_in_net,
      en(0) => convert1_dout_net,
      rst => "0",
      q => register1_q_net
    );

  register12: entity warp_per_block_calc_lib.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d(0) => relational_op_net,
      en => "1",
      rst => "0",
      q(0) => data_valid_out_net
    );

  register2: entity warp_per_block_calc_lib.xlregister
    generic map (
      d_width => 6,
      init_value => b"000000"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d => mux_y_net,
      en(0) => relational_op_net,
      rst => "0",
      q => warps_per_block_out_net
    );

  register3: entity warp_per_block_calc_lib.xlregister
    generic map (
      d_width => 6,
      init_value => b"000000"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d => warp_size_in_net,
      en(0) => convert1_dout_net,
      rst => "0",
      q => register3_q_net
    );

  register7: entity warp_per_block_calc_lib.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d(0) => convert1_dout_net,
      en(0) => logical_y_net,
      rst => "0",
      q(0) => register7_q_net
    );

  relational: entity warp_per_block_calc_lib.relational_54048c8b02
    port map (
      a => constant2_op_net,
      b => counter3_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational_op_net
    );

  relational1: entity warp_per_block_calc_lib.relational_4eca908438
    port map (
      a => divider_generator_3_0_fractional_net,
      b(0) => constant1_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => relational1_op_net
    );

end structural;
