--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2012 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file addsb_11_0_f45daeb7eb283db0.vhd when simulating
-- the core, addsb_11_0_f45daeb7eb283db0. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY addsb_11_0_f45daeb7eb283db0 IS
  PORT (
    a : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(32 DOWNTO 0)
  );
END addsb_11_0_f45daeb7eb283db0;

ARCHITECTURE addsb_11_0_f45daeb7eb283db0_a OF addsb_11_0_f45daeb7eb283db0 IS
-- synthesis translate_off
COMPONENT wrapped_addsb_11_0_f45daeb7eb283db0
  PORT (
    a : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    s : OUT STD_LOGIC_VECTOR(32 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_addsb_11_0_f45daeb7eb283db0 USE ENTITY XilinxCoreLib.c_addsub_v11_0(behavioral)
    GENERIC MAP (
      c_a_type => 1,
      c_a_width => 33,
      c_add_mode => 0,
      c_ainit_val => "0",
      c_b_constant => 0,
      c_b_type => 1,
      c_b_value => "000000000000000000000000000000000",
      c_b_width => 33,
      c_borrow_low => 1,
      c_bypass_low => 0,
      c_ce_overrides_bypass => 1,
      c_ce_overrides_sclr => 0,
      c_has_bypass => 0,
      c_has_c_in => 0,
      c_has_c_out => 0,
      c_has_ce => 0,
      c_has_sclr => 0,
      c_has_sinit => 0,
      c_has_sset => 0,
      c_implementation => 0,
      c_latency => 0,
      c_out_width => 33,
      c_sclr_overrides_sset => 0,
      c_sinit_val => "0",
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_addsb_11_0_f45daeb7eb283db0
  PORT MAP (
    a => a,
    b => b,
    s => s
  );
-- synthesis translate_on

END addsb_11_0_f45daeb7eb283db0_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2012 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file cntr_11_0_e7514e290b172ea1.vhd when simulating
-- the core, cntr_11_0_e7514e290b172ea1. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY cntr_11_0_e7514e290b172ea1 IS
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END cntr_11_0_e7514e290b172ea1;

ARCHITECTURE cntr_11_0_e7514e290b172ea1_a OF cntr_11_0_e7514e290b172ea1 IS
-- synthesis translate_off
COMPONENT wrapped_cntr_11_0_e7514e290b172ea1
  PORT (
    clk : IN STD_LOGIC;
    ce : IN STD_LOGIC;
    sinit : IN STD_LOGIC;
    q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_cntr_11_0_e7514e290b172ea1 USE ENTITY XilinxCoreLib.c_counter_binary_v11_0(behavioral)
    GENERIC MAP (
      c_ainit_val => "0",
      c_ce_overrides_sync => 0,
      c_count_by => "1",
      c_count_mode => 0,
      c_count_to => "1",
      c_fb_latency => 0,
      c_has_ce => 1,
      c_has_load => 0,
      c_has_sclr => 0,
      c_has_sinit => 1,
      c_has_sset => 0,
      c_has_thresh0 => 0,
      c_implementation => 0,
      c_latency => 1,
      c_load_low => 0,
      c_restrict_count => 0,
      c_sclr_overrides_sset => 1,
      c_sinit_val => "0",
      c_thresh0_value => "1",
      c_verbosity => 0,
      c_width => 8,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_cntr_11_0_e7514e290b172ea1
  PORT MAP (
    clk => clk,
    ce => ce,
    sinit => sinit,
    q => q
  );
-- synthesis translate_on

END cntr_11_0_e7514e290b172ea1_a;
--------------------------------------------------------------------------------
-- Copyright (c) 1995-2011 Xilinx, Inc.  All rights reserved.
--------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version: O.61xd
--  \   \         Application: netgen
--  /   /         Filename: dv_gn_v3_0_26253f791d7c00ab.vhd
-- /___/   /\     Timestamp: Mon Jul 23 19:55:10 2012
-- \   \  /  \ 
--  \___\/\___\
--             
-- Command	: -intstyle ise -w -sim -ofmt vhdl ./tmp/_cg/dv_gn_v3_0_26253f791d7c00ab.ngc ./tmp/_cg/dv_gn_v3_0_26253f791d7c00ab.vhd 
-- Device	: 6vcx75tff484-2
-- Input file	: ./tmp/_cg/dv_gn_v3_0_26253f791d7c00ab.ngc
-- Output file	: ./tmp/_cg/dv_gn_v3_0_26253f791d7c00ab.vhd
-- # of Entities	: 1
-- Design Name	: dv_gn_v3_0_26253f791d7c00ab
-- Xilinx	: c:\xilinx\13.2\ise_ds\ise\
--             
-- Purpose:    
--     This VHDL netlist is a verification model and uses simulation 
--     primitives which may not represent the true implementation of the 
--     device, however the netlist is functionally correct and should not 
--     be modified. This file cannot be synthesized and should only be used 
--     with supported simulation tools.
--             
-- Reference:  
--     Command Line Tools User Guide, Chapter 23
--     Synthesis and Simulation Design Guide, Chapter 6
--             
--------------------------------------------------------------------------------


-- synthesis translate_off
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;
use UNISIM.VPKG.ALL;

entity dv_gn_v3_0_26253f791d7c00ab is
  port (
    ce : in STD_LOGIC := 'X'; 
    rfd : out STD_LOGIC; 
    clk : in STD_LOGIC := 'X'; 
    dividend : in STD_LOGIC_VECTOR ( 5 downto 0 ); 
    quotient : out STD_LOGIC_VECTOR ( 5 downto 0 ); 
    divisor : in STD_LOGIC_VECTOR ( 7 downto 0 ); 
    fractional : out STD_LOGIC_VECTOR ( 7 downto 0 ) 
  );
end dv_gn_v3_0_26253f791d7c00ab;

architecture STRUCTURE of dv_gn_v3_0_26253f791d7c00ab is
  signal NlwRenamedSig_OI_rfd : STD_LOGIC; 
  signal blk00000003_sig00000188 : STD_LOGIC; 
  signal blk00000003_sig00000187 : STD_LOGIC; 
  signal blk00000003_sig00000186 : STD_LOGIC; 
  signal blk00000003_sig00000185 : STD_LOGIC; 
  signal blk00000003_sig00000184 : STD_LOGIC; 
  signal blk00000003_sig00000183 : STD_LOGIC; 
  signal blk00000003_sig00000182 : STD_LOGIC; 
  signal blk00000003_sig00000181 : STD_LOGIC; 
  signal blk00000003_sig00000180 : STD_LOGIC; 
  signal blk00000003_sig0000017f : STD_LOGIC; 
  signal blk00000003_sig0000017e : STD_LOGIC; 
  signal blk00000003_sig0000017d : STD_LOGIC; 
  signal blk00000003_sig0000017c : STD_LOGIC; 
  signal blk00000003_sig0000017b : STD_LOGIC; 
  signal blk00000003_sig0000017a : STD_LOGIC; 
  signal blk00000003_sig00000179 : STD_LOGIC; 
  signal blk00000003_sig00000178 : STD_LOGIC; 
  signal blk00000003_sig00000177 : STD_LOGIC; 
  signal blk00000003_sig00000176 : STD_LOGIC; 
  signal blk00000003_sig00000175 : STD_LOGIC; 
  signal blk00000003_sig00000174 : STD_LOGIC; 
  signal blk00000003_sig00000173 : STD_LOGIC; 
  signal blk00000003_sig00000172 : STD_LOGIC; 
  signal blk00000003_sig00000171 : STD_LOGIC; 
  signal blk00000003_sig00000170 : STD_LOGIC; 
  signal blk00000003_sig0000016f : STD_LOGIC; 
  signal blk00000003_sig0000016e : STD_LOGIC; 
  signal blk00000003_sig0000016d : STD_LOGIC; 
  signal blk00000003_sig0000016c : STD_LOGIC; 
  signal blk00000003_sig0000016b : STD_LOGIC; 
  signal blk00000003_sig0000016a : STD_LOGIC; 
  signal blk00000003_sig00000169 : STD_LOGIC; 
  signal blk00000003_sig00000168 : STD_LOGIC; 
  signal blk00000003_sig00000167 : STD_LOGIC; 
  signal blk00000003_sig00000166 : STD_LOGIC; 
  signal blk00000003_sig00000165 : STD_LOGIC; 
  signal blk00000003_sig00000164 : STD_LOGIC; 
  signal blk00000003_sig00000163 : STD_LOGIC; 
  signal blk00000003_sig00000162 : STD_LOGIC; 
  signal blk00000003_sig00000161 : STD_LOGIC; 
  signal blk00000003_sig00000160 : STD_LOGIC; 
  signal blk00000003_sig0000015f : STD_LOGIC; 
  signal blk00000003_sig0000015e : STD_LOGIC; 
  signal blk00000003_sig0000015d : STD_LOGIC; 
  signal blk00000003_sig0000015c : STD_LOGIC; 
  signal blk00000003_sig0000015b : STD_LOGIC; 
  signal blk00000003_sig0000015a : STD_LOGIC; 
  signal blk00000003_sig00000159 : STD_LOGIC; 
  signal blk00000003_sig00000158 : STD_LOGIC; 
  signal blk00000003_sig00000157 : STD_LOGIC; 
  signal blk00000003_sig00000156 : STD_LOGIC; 
  signal blk00000003_sig00000155 : STD_LOGIC; 
  signal blk00000003_sig00000154 : STD_LOGIC; 
  signal blk00000003_sig00000153 : STD_LOGIC; 
  signal blk00000003_sig00000152 : STD_LOGIC; 
  signal blk00000003_sig00000151 : STD_LOGIC; 
  signal blk00000003_sig00000150 : STD_LOGIC; 
  signal blk00000003_sig0000014f : STD_LOGIC; 
  signal blk00000003_sig0000014e : STD_LOGIC; 
  signal blk00000003_sig0000014d : STD_LOGIC; 
  signal blk00000003_sig0000014c : STD_LOGIC; 
  signal blk00000003_sig0000014b : STD_LOGIC; 
  signal blk00000003_sig0000014a : STD_LOGIC; 
  signal blk00000003_sig00000149 : STD_LOGIC; 
  signal blk00000003_sig00000148 : STD_LOGIC; 
  signal blk00000003_sig00000147 : STD_LOGIC; 
  signal blk00000003_sig00000146 : STD_LOGIC; 
  signal blk00000003_sig00000145 : STD_LOGIC; 
  signal blk00000003_sig00000144 : STD_LOGIC; 
  signal blk00000003_sig00000143 : STD_LOGIC; 
  signal blk00000003_sig00000142 : STD_LOGIC; 
  signal blk00000003_sig00000141 : STD_LOGIC; 
  signal blk00000003_sig00000140 : STD_LOGIC; 
  signal blk00000003_sig0000013f : STD_LOGIC; 
  signal blk00000003_sig0000013e : STD_LOGIC; 
  signal blk00000003_sig0000013d : STD_LOGIC; 
  signal blk00000003_sig0000013c : STD_LOGIC; 
  signal blk00000003_sig0000013b : STD_LOGIC; 
  signal blk00000003_sig0000013a : STD_LOGIC; 
  signal blk00000003_sig00000139 : STD_LOGIC; 
  signal blk00000003_sig00000138 : STD_LOGIC; 
  signal blk00000003_sig00000137 : STD_LOGIC; 
  signal blk00000003_sig00000136 : STD_LOGIC; 
  signal blk00000003_sig00000135 : STD_LOGIC; 
  signal blk00000003_sig00000134 : STD_LOGIC; 
  signal blk00000003_sig00000133 : STD_LOGIC; 
  signal blk00000003_sig00000132 : STD_LOGIC; 
  signal blk00000003_sig00000131 : STD_LOGIC; 
  signal blk00000003_sig00000130 : STD_LOGIC; 
  signal blk00000003_sig0000012f : STD_LOGIC; 
  signal blk00000003_sig0000012e : STD_LOGIC; 
  signal blk00000003_sig0000012d : STD_LOGIC; 
  signal blk00000003_sig0000012c : STD_LOGIC; 
  signal blk00000003_sig0000012b : STD_LOGIC; 
  signal blk00000003_sig0000012a : STD_LOGIC; 
  signal blk00000003_sig00000129 : STD_LOGIC; 
  signal blk00000003_sig00000128 : STD_LOGIC; 
  signal blk00000003_sig00000127 : STD_LOGIC; 
  signal blk00000003_sig00000126 : STD_LOGIC; 
  signal blk00000003_sig00000125 : STD_LOGIC; 
  signal blk00000003_sig00000124 : STD_LOGIC; 
  signal blk00000003_sig00000123 : STD_LOGIC; 
  signal blk00000003_sig00000122 : STD_LOGIC; 
  signal blk00000003_sig00000121 : STD_LOGIC; 
  signal blk00000003_sig00000120 : STD_LOGIC; 
  signal blk00000003_sig0000011f : STD_LOGIC; 
  signal blk00000003_sig0000011e : STD_LOGIC; 
  signal blk00000003_sig0000011d : STD_LOGIC; 
  signal blk00000003_sig0000011c : STD_LOGIC; 
  signal blk00000003_sig0000011b : STD_LOGIC; 
  signal blk00000003_sig0000011a : STD_LOGIC; 
  signal blk00000003_sig00000119 : STD_LOGIC; 
  signal blk00000003_sig00000118 : STD_LOGIC; 
  signal blk00000003_sig00000117 : STD_LOGIC; 
  signal blk00000003_sig00000116 : STD_LOGIC; 
  signal blk00000003_sig00000115 : STD_LOGIC; 
  signal blk00000003_sig00000114 : STD_LOGIC; 
  signal blk00000003_sig00000113 : STD_LOGIC; 
  signal blk00000003_sig00000112 : STD_LOGIC; 
  signal blk00000003_sig00000111 : STD_LOGIC; 
  signal blk00000003_sig00000110 : STD_LOGIC; 
  signal blk00000003_sig0000010f : STD_LOGIC; 
  signal blk00000003_sig0000010e : STD_LOGIC; 
  signal blk00000003_sig0000010d : STD_LOGIC; 
  signal blk00000003_sig0000010c : STD_LOGIC; 
  signal blk00000003_sig0000010b : STD_LOGIC; 
  signal blk00000003_sig0000010a : STD_LOGIC; 
  signal blk00000003_sig00000109 : STD_LOGIC; 
  signal blk00000003_sig00000108 : STD_LOGIC; 
  signal blk00000003_sig00000107 : STD_LOGIC; 
  signal blk00000003_sig00000106 : STD_LOGIC; 
  signal blk00000003_sig00000105 : STD_LOGIC; 
  signal blk00000003_sig00000104 : STD_LOGIC; 
  signal blk00000003_sig00000103 : STD_LOGIC; 
  signal blk00000003_sig00000102 : STD_LOGIC; 
  signal blk00000003_sig00000101 : STD_LOGIC; 
  signal blk00000003_sig00000100 : STD_LOGIC; 
  signal blk00000003_sig000000ff : STD_LOGIC; 
  signal blk00000003_sig000000fe : STD_LOGIC; 
  signal blk00000003_sig000000fd : STD_LOGIC; 
  signal blk00000003_sig000000fc : STD_LOGIC; 
  signal blk00000003_sig000000fb : STD_LOGIC; 
  signal blk00000003_sig000000fa : STD_LOGIC; 
  signal blk00000003_sig000000f9 : STD_LOGIC; 
  signal blk00000003_sig000000f8 : STD_LOGIC; 
  signal blk00000003_sig000000f7 : STD_LOGIC; 
  signal blk00000003_sig000000f6 : STD_LOGIC; 
  signal blk00000003_sig000000f5 : STD_LOGIC; 
  signal blk00000003_sig000000f4 : STD_LOGIC; 
  signal blk00000003_sig000000f3 : STD_LOGIC; 
  signal blk00000003_sig000000f2 : STD_LOGIC; 
  signal blk00000003_sig000000f1 : STD_LOGIC; 
  signal blk00000003_sig000000f0 : STD_LOGIC; 
  signal blk00000003_sig000000ef : STD_LOGIC; 
  signal blk00000003_sig000000ee : STD_LOGIC; 
  signal blk00000003_sig000000ed : STD_LOGIC; 
  signal blk00000003_sig000000ec : STD_LOGIC; 
  signal blk00000003_sig000000eb : STD_LOGIC; 
  signal blk00000003_sig000000ea : STD_LOGIC; 
  signal blk00000003_sig000000e9 : STD_LOGIC; 
  signal blk00000003_sig000000e8 : STD_LOGIC; 
  signal blk00000003_sig000000e7 : STD_LOGIC; 
  signal blk00000003_sig000000e6 : STD_LOGIC; 
  signal blk00000003_sig000000e5 : STD_LOGIC; 
  signal blk00000003_sig000000e4 : STD_LOGIC; 
  signal blk00000003_sig000000e3 : STD_LOGIC; 
  signal blk00000003_sig000000e2 : STD_LOGIC; 
  signal blk00000003_sig000000e1 : STD_LOGIC; 
  signal blk00000003_sig000000e0 : STD_LOGIC; 
  signal blk00000003_sig000000df : STD_LOGIC; 
  signal blk00000003_sig000000de : STD_LOGIC; 
  signal blk00000003_sig000000dd : STD_LOGIC; 
  signal blk00000003_sig000000dc : STD_LOGIC; 
  signal blk00000003_sig000000db : STD_LOGIC; 
  signal blk00000003_sig000000da : STD_LOGIC; 
  signal blk00000003_sig000000d9 : STD_LOGIC; 
  signal blk00000003_sig000000d8 : STD_LOGIC; 
  signal blk00000003_sig000000d7 : STD_LOGIC; 
  signal blk00000003_sig000000d6 : STD_LOGIC; 
  signal blk00000003_sig000000d5 : STD_LOGIC; 
  signal blk00000003_sig000000d4 : STD_LOGIC; 
  signal blk00000003_sig000000d3 : STD_LOGIC; 
  signal blk00000003_sig000000d2 : STD_LOGIC; 
  signal blk00000003_sig000000d1 : STD_LOGIC; 
  signal blk00000003_sig000000d0 : STD_LOGIC; 
  signal blk00000003_sig000000cf : STD_LOGIC; 
  signal blk00000003_sig000000ce : STD_LOGIC; 
  signal blk00000003_sig000000cd : STD_LOGIC; 
  signal blk00000003_sig000000cc : STD_LOGIC; 
  signal blk00000003_sig000000cb : STD_LOGIC; 
  signal blk00000003_sig000000ca : STD_LOGIC; 
  signal blk00000003_sig000000c9 : STD_LOGIC; 
  signal blk00000003_sig000000c8 : STD_LOGIC; 
  signal blk00000003_sig000000c7 : STD_LOGIC; 
  signal blk00000003_sig000000c6 : STD_LOGIC; 
  signal blk00000003_sig000000c5 : STD_LOGIC; 
  signal blk00000003_sig000000c4 : STD_LOGIC; 
  signal blk00000003_sig000000c3 : STD_LOGIC; 
  signal blk00000003_sig000000c2 : STD_LOGIC; 
  signal blk00000003_sig000000c1 : STD_LOGIC; 
  signal blk00000003_sig000000c0 : STD_LOGIC; 
  signal blk00000003_sig000000bf : STD_LOGIC; 
  signal blk00000003_sig000000be : STD_LOGIC; 
  signal blk00000003_sig000000bd : STD_LOGIC; 
  signal blk00000003_sig000000bc : STD_LOGIC; 
  signal blk00000003_sig000000bb : STD_LOGIC; 
  signal blk00000003_sig000000ba : STD_LOGIC; 
  signal blk00000003_sig000000b9 : STD_LOGIC; 
  signal blk00000003_sig000000b8 : STD_LOGIC; 
  signal blk00000003_sig000000b7 : STD_LOGIC; 
  signal blk00000003_sig000000b6 : STD_LOGIC; 
  signal blk00000003_sig000000b5 : STD_LOGIC; 
  signal blk00000003_sig000000b4 : STD_LOGIC; 
  signal blk00000003_sig000000b3 : STD_LOGIC; 
  signal blk00000003_sig000000b2 : STD_LOGIC; 
  signal blk00000003_sig000000b1 : STD_LOGIC; 
  signal blk00000003_sig000000b0 : STD_LOGIC; 
  signal blk00000003_sig000000af : STD_LOGIC; 
  signal blk00000003_sig000000ae : STD_LOGIC; 
  signal blk00000003_sig000000ad : STD_LOGIC; 
  signal blk00000003_sig000000ac : STD_LOGIC; 
  signal blk00000003_sig000000ab : STD_LOGIC; 
  signal blk00000003_sig000000aa : STD_LOGIC; 
  signal blk00000003_sig000000a9 : STD_LOGIC; 
  signal blk00000003_sig000000a8 : STD_LOGIC; 
  signal blk00000003_sig000000a7 : STD_LOGIC; 
  signal blk00000003_sig000000a6 : STD_LOGIC; 
  signal blk00000003_sig000000a5 : STD_LOGIC; 
  signal blk00000003_sig000000a4 : STD_LOGIC; 
  signal blk00000003_sig000000a3 : STD_LOGIC; 
  signal blk00000003_sig000000a2 : STD_LOGIC; 
  signal blk00000003_sig000000a1 : STD_LOGIC; 
  signal blk00000003_sig000000a0 : STD_LOGIC; 
  signal blk00000003_sig0000009f : STD_LOGIC; 
  signal blk00000003_sig0000009e : STD_LOGIC; 
  signal blk00000003_sig0000009d : STD_LOGIC; 
  signal blk00000003_sig0000009c : STD_LOGIC; 
  signal blk00000003_sig0000009b : STD_LOGIC; 
  signal blk00000003_sig0000009a : STD_LOGIC; 
  signal blk00000003_sig00000099 : STD_LOGIC; 
  signal blk00000003_sig00000098 : STD_LOGIC; 
  signal blk00000003_sig00000097 : STD_LOGIC; 
  signal blk00000003_sig00000096 : STD_LOGIC; 
  signal blk00000003_sig00000095 : STD_LOGIC; 
  signal blk00000003_sig00000094 : STD_LOGIC; 
  signal blk00000003_sig00000093 : STD_LOGIC; 
  signal blk00000003_sig00000092 : STD_LOGIC; 
  signal blk00000003_sig00000091 : STD_LOGIC; 
  signal blk00000003_sig00000090 : STD_LOGIC; 
  signal blk00000003_sig0000008f : STD_LOGIC; 
  signal blk00000003_sig0000008e : STD_LOGIC; 
  signal blk00000003_sig0000008d : STD_LOGIC; 
  signal blk00000003_sig0000008c : STD_LOGIC; 
  signal blk00000003_sig0000008b : STD_LOGIC; 
  signal blk00000003_sig0000008a : STD_LOGIC; 
  signal blk00000003_sig00000089 : STD_LOGIC; 
  signal blk00000003_sig00000088 : STD_LOGIC; 
  signal blk00000003_sig00000087 : STD_LOGIC; 
  signal blk00000003_sig00000086 : STD_LOGIC; 
  signal blk00000003_sig00000085 : STD_LOGIC; 
  signal blk00000003_sig00000084 : STD_LOGIC; 
  signal blk00000003_sig00000083 : STD_LOGIC; 
  signal blk00000003_sig00000082 : STD_LOGIC; 
  signal blk00000003_sig00000081 : STD_LOGIC; 
  signal blk00000003_sig00000080 : STD_LOGIC; 
  signal blk00000003_sig0000007f : STD_LOGIC; 
  signal blk00000003_sig0000007e : STD_LOGIC; 
  signal blk00000003_sig0000007d : STD_LOGIC; 
  signal blk00000003_sig0000007c : STD_LOGIC; 
  signal blk00000003_sig0000007b : STD_LOGIC; 
  signal blk00000003_sig0000007a : STD_LOGIC; 
  signal blk00000003_sig00000079 : STD_LOGIC; 
  signal blk00000003_sig00000078 : STD_LOGIC; 
  signal blk00000003_sig00000077 : STD_LOGIC; 
  signal blk00000003_sig00000076 : STD_LOGIC; 
  signal blk00000003_sig00000075 : STD_LOGIC; 
  signal blk00000003_sig00000074 : STD_LOGIC; 
  signal blk00000003_sig00000073 : STD_LOGIC; 
  signal blk00000003_sig00000072 : STD_LOGIC; 
  signal blk00000003_sig00000071 : STD_LOGIC; 
  signal blk00000003_sig00000070 : STD_LOGIC; 
  signal blk00000003_sig0000006f : STD_LOGIC; 
  signal blk00000003_sig0000006e : STD_LOGIC; 
  signal blk00000003_sig0000006d : STD_LOGIC; 
  signal blk00000003_sig0000006c : STD_LOGIC; 
  signal blk00000003_sig0000006b : STD_LOGIC; 
  signal blk00000003_sig0000006a : STD_LOGIC; 
  signal blk00000003_sig00000069 : STD_LOGIC; 
  signal blk00000003_sig00000068 : STD_LOGIC; 
  signal blk00000003_sig00000067 : STD_LOGIC; 
  signal blk00000003_sig00000066 : STD_LOGIC; 
  signal blk00000003_sig00000065 : STD_LOGIC; 
  signal blk00000003_sig00000064 : STD_LOGIC; 
  signal blk00000003_sig00000063 : STD_LOGIC; 
  signal blk00000003_sig00000062 : STD_LOGIC; 
  signal blk00000003_sig00000061 : STD_LOGIC; 
  signal blk00000003_sig00000060 : STD_LOGIC; 
  signal blk00000003_sig0000005f : STD_LOGIC; 
  signal blk00000003_sig0000005e : STD_LOGIC; 
  signal blk00000003_sig0000005d : STD_LOGIC; 
  signal blk00000003_sig0000005c : STD_LOGIC; 
  signal blk00000003_sig0000005b : STD_LOGIC; 
  signal blk00000003_sig0000005a : STD_LOGIC; 
  signal blk00000003_sig00000059 : STD_LOGIC; 
  signal blk00000003_sig00000058 : STD_LOGIC; 
  signal blk00000003_sig00000057 : STD_LOGIC; 
  signal blk00000003_sig00000056 : STD_LOGIC; 
  signal blk00000003_sig00000055 : STD_LOGIC; 
  signal blk00000003_sig00000054 : STD_LOGIC; 
  signal blk00000003_sig00000053 : STD_LOGIC; 
  signal blk00000003_sig00000052 : STD_LOGIC; 
  signal blk00000003_sig00000051 : STD_LOGIC; 
  signal blk00000003_sig00000050 : STD_LOGIC; 
  signal blk00000003_sig0000004f : STD_LOGIC; 
  signal blk00000003_sig0000004e : STD_LOGIC; 
  signal blk00000003_sig0000004d : STD_LOGIC; 
  signal blk00000003_sig0000004c : STD_LOGIC; 
  signal blk00000003_sig0000004b : STD_LOGIC; 
  signal blk00000003_sig0000004a : STD_LOGIC; 
  signal blk00000003_sig00000049 : STD_LOGIC; 
  signal blk00000003_sig00000048 : STD_LOGIC; 
  signal blk00000003_sig00000047 : STD_LOGIC; 
  signal blk00000003_sig00000046 : STD_LOGIC; 
  signal blk00000003_sig00000045 : STD_LOGIC; 
  signal blk00000003_sig00000044 : STD_LOGIC; 
  signal blk00000003_sig00000043 : STD_LOGIC; 
  signal blk00000003_sig00000042 : STD_LOGIC; 
  signal blk00000003_sig00000041 : STD_LOGIC; 
  signal blk00000003_sig00000040 : STD_LOGIC; 
  signal blk00000003_sig0000003f : STD_LOGIC; 
  signal blk00000003_sig0000003e : STD_LOGIC; 
  signal blk00000003_sig0000003d : STD_LOGIC; 
  signal blk00000003_sig0000003c : STD_LOGIC; 
  signal blk00000003_sig0000003b : STD_LOGIC; 
  signal blk00000003_sig0000003a : STD_LOGIC; 
  signal blk00000003_sig00000039 : STD_LOGIC; 
  signal blk00000003_sig00000038 : STD_LOGIC; 
  signal blk00000003_sig00000037 : STD_LOGIC; 
  signal blk00000003_sig00000036 : STD_LOGIC; 
  signal blk00000003_sig00000035 : STD_LOGIC; 
  signal blk00000003_sig00000034 : STD_LOGIC; 
  signal blk00000003_sig00000033 : STD_LOGIC; 
  signal blk00000003_sig00000032 : STD_LOGIC; 
  signal blk00000003_sig00000031 : STD_LOGIC; 
  signal blk00000003_sig00000030 : STD_LOGIC; 
  signal blk00000003_sig0000002f : STD_LOGIC; 
  signal blk00000003_sig0000002e : STD_LOGIC; 
  signal blk00000003_sig0000002d : STD_LOGIC; 
  signal blk00000003_sig0000002c : STD_LOGIC; 
  signal blk00000003_sig0000002b : STD_LOGIC; 
  signal blk00000003_sig0000002a : STD_LOGIC; 
  signal blk00000003_sig00000029 : STD_LOGIC; 
  signal blk00000003_sig00000028 : STD_LOGIC; 
  signal blk00000003_sig00000027 : STD_LOGIC; 
  signal blk00000003_sig00000026 : STD_LOGIC; 
  signal blk00000003_sig00000025 : STD_LOGIC; 
  signal blk00000003_sig00000024 : STD_LOGIC; 
  signal blk00000003_sig00000023 : STD_LOGIC; 
  signal blk00000003_sig00000022 : STD_LOGIC; 
  signal blk00000003_sig00000021 : STD_LOGIC; 
  signal blk00000003_sig0000001f : STD_LOGIC; 
  signal NLW_blk00000001_P_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000002_G_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000003_blk00000068_O_UNCONNECTED : STD_LOGIC; 
begin
  rfd <= NlwRenamedSig_OI_rfd;
  blk00000001 : VCC
    port map (
      P => NLW_blk00000001_P_UNCONNECTED
    );
  blk00000002 : GND
    port map (
      G => NLW_blk00000002_G_UNCONNECTED
    );
  blk00000003_blk0000017c : INV
    port map (
      I => blk00000003_sig00000080,
      O => blk00000003_sig0000008a
    );
  blk00000003_blk0000017b : INV
    port map (
      I => blk00000003_sig00000081,
      O => blk00000003_sig0000008d
    );
  blk00000003_blk0000017a : INV
    port map (
      I => blk00000003_sig00000082,
      O => blk00000003_sig00000090
    );
  blk00000003_blk00000179 : INV
    port map (
      I => blk00000003_sig00000083,
      O => blk00000003_sig00000093
    );
  blk00000003_blk00000178 : INV
    port map (
      I => blk00000003_sig00000084,
      O => blk00000003_sig00000096
    );
  blk00000003_blk00000177 : INV
    port map (
      I => blk00000003_sig00000085,
      O => blk00000003_sig00000099
    );
  blk00000003_blk00000176 : INV
    port map (
      I => blk00000003_sig00000086,
      O => blk00000003_sig0000009c
    );
  blk00000003_blk00000175 : INV
    port map (
      I => blk00000003_sig0000002a,
      O => blk00000003_sig0000004f
    );
  blk00000003_blk00000174 : INV
    port map (
      I => blk00000003_sig00000028,
      O => blk00000003_sig0000004e
    );
  blk00000003_blk00000173 : INV
    port map (
      I => blk00000003_sig00000026,
      O => blk00000003_sig0000004d
    );
  blk00000003_blk00000172 : INV
    port map (
      I => blk00000003_sig00000024,
      O => blk00000003_sig0000004c
    );
  blk00000003_blk00000171 : INV
    port map (
      I => blk00000003_sig00000022,
      O => blk00000003_sig0000004b
    );
  blk00000003_blk00000170 : INV
    port map (
      I => blk00000003_sig00000021,
      O => blk00000003_sig00000157
    );
  blk00000003_blk0000016f : INV
    port map (
      I => blk00000003_sig0000002b,
      O => blk00000003_sig00000132
    );
  blk00000003_blk0000016e : INV
    port map (
      I => blk00000003_sig00000033,
      O => blk00000003_sig0000010d
    );
  blk00000003_blk0000016d : INV
    port map (
      I => blk00000003_sig0000003a,
      O => blk00000003_sig000000e8
    );
  blk00000003_blk0000016c : INV
    port map (
      I => blk00000003_sig00000041,
      O => blk00000003_sig000000c3
    );
  blk00000003_blk0000016b : LUT1
    generic map(
      INIT => X"1"
    )
    port map (
      I0 => blk00000003_sig000000a1,
      O => blk00000003_sig00000041
    );
  blk00000003_blk0000016a : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig0000015c,
      I1 => blk00000003_sig00000051,
      I2 => blk00000003_sig0000015b,
      O => blk00000003_sig00000165
    );
  blk00000003_blk00000169 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig0000015d,
      I1 => blk00000003_sig00000053,
      I2 => blk00000003_sig0000015b,
      O => blk00000003_sig00000168
    );
  blk00000003_blk00000168 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig0000015e,
      I1 => blk00000003_sig00000055,
      I2 => blk00000003_sig0000015b,
      O => blk00000003_sig0000016b
    );
  blk00000003_blk00000167 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig0000015f,
      I1 => blk00000003_sig00000057,
      I2 => blk00000003_sig0000015b,
      O => blk00000003_sig0000016e
    );
  blk00000003_blk00000166 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000160,
      I1 => blk00000003_sig00000059,
      I2 => blk00000003_sig0000015b,
      O => blk00000003_sig00000171
    );
  blk00000003_blk00000165 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000161,
      I1 => blk00000003_sig0000005b,
      I2 => blk00000003_sig0000015b,
      O => blk00000003_sig00000174
    );
  blk00000003_blk00000164 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000162,
      I1 => blk00000003_sig0000005d,
      I2 => blk00000003_sig0000015b,
      O => blk00000003_sig00000177
    );
  blk00000003_blk00000163 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000163,
      I1 => blk00000003_sig0000005f,
      I2 => blk00000003_sig0000015b,
      O => blk00000003_sig00000184
    );
  blk00000003_blk00000162 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000155,
      I1 => blk00000003_sig00000021,
      O => blk00000003_sig00000137
    );
  blk00000003_blk00000161 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000014e,
      I1 => blk00000003_sig00000050,
      I2 => blk00000003_sig00000021,
      O => blk00000003_sig0000013a
    );
  blk00000003_blk00000160 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000014f,
      I1 => blk00000003_sig00000052,
      I2 => blk00000003_sig00000021,
      O => blk00000003_sig0000013d
    );
  blk00000003_blk0000015f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000150,
      I1 => blk00000003_sig00000054,
      I2 => blk00000003_sig00000021,
      O => blk00000003_sig00000140
    );
  blk00000003_blk0000015e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000151,
      I1 => blk00000003_sig00000056,
      I2 => blk00000003_sig00000021,
      O => blk00000003_sig00000143
    );
  blk00000003_blk0000015d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000152,
      I1 => blk00000003_sig00000058,
      I2 => blk00000003_sig00000021,
      O => blk00000003_sig00000146
    );
  blk00000003_blk0000015c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000153,
      I1 => blk00000003_sig0000005a,
      I2 => blk00000003_sig00000021,
      O => blk00000003_sig00000149
    );
  blk00000003_blk0000015b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000154,
      I1 => blk00000003_sig0000005c,
      I2 => blk00000003_sig00000021,
      O => blk00000003_sig0000014c
    );
  blk00000003_blk0000015a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000048,
      I1 => blk00000003_sig0000005e,
      I2 => blk00000003_sig00000021,
      O => blk00000003_sig00000158
    );
  blk00000003_blk00000159 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000130,
      I1 => blk00000003_sig0000002b,
      O => blk00000003_sig00000112
    );
  blk00000003_blk00000158 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000129,
      I1 => blk00000003_sig00000060,
      I2 => blk00000003_sig0000002b,
      O => blk00000003_sig00000115
    );
  blk00000003_blk00000157 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000012a,
      I1 => blk00000003_sig00000061,
      I2 => blk00000003_sig0000002b,
      O => blk00000003_sig00000118
    );
  blk00000003_blk00000156 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000012b,
      I1 => blk00000003_sig00000062,
      I2 => blk00000003_sig0000002b,
      O => blk00000003_sig0000011b
    );
  blk00000003_blk00000155 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000012c,
      I1 => blk00000003_sig00000063,
      I2 => blk00000003_sig0000002b,
      O => blk00000003_sig0000011e
    );
  blk00000003_blk00000154 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000012d,
      I1 => blk00000003_sig00000064,
      I2 => blk00000003_sig0000002b,
      O => blk00000003_sig00000121
    );
  blk00000003_blk00000153 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000012e,
      I1 => blk00000003_sig00000065,
      I2 => blk00000003_sig0000002b,
      O => blk00000003_sig00000124
    );
  blk00000003_blk00000152 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000012f,
      I1 => blk00000003_sig00000066,
      I2 => blk00000003_sig0000002b,
      O => blk00000003_sig00000127
    );
  blk00000003_blk00000151 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000032,
      I1 => blk00000003_sig00000067,
      I2 => blk00000003_sig0000002b,
      O => blk00000003_sig00000133
    );
  blk00000003_blk00000150 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000010b,
      I1 => blk00000003_sig00000033,
      O => blk00000003_sig000000ed
    );
  blk00000003_blk0000014f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000104,
      I1 => blk00000003_sig00000068,
      I2 => blk00000003_sig00000033,
      O => blk00000003_sig000000f0
    );
  blk00000003_blk0000014e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000105,
      I1 => blk00000003_sig00000069,
      I2 => blk00000003_sig00000033,
      O => blk00000003_sig000000f3
    );
  blk00000003_blk0000014d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000106,
      I1 => blk00000003_sig0000006a,
      I2 => blk00000003_sig00000033,
      O => blk00000003_sig000000f6
    );
  blk00000003_blk0000014c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000107,
      I1 => blk00000003_sig0000006b,
      I2 => blk00000003_sig00000033,
      O => blk00000003_sig000000f9
    );
  blk00000003_blk0000014b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000108,
      I1 => blk00000003_sig0000006c,
      I2 => blk00000003_sig00000033,
      O => blk00000003_sig000000fc
    );
  blk00000003_blk0000014a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000109,
      I1 => blk00000003_sig0000006d,
      I2 => blk00000003_sig00000033,
      O => blk00000003_sig000000ff
    );
  blk00000003_blk00000149 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000010a,
      I1 => blk00000003_sig0000006e,
      I2 => blk00000003_sig00000033,
      O => blk00000003_sig00000102
    );
  blk00000003_blk00000148 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000039,
      I1 => blk00000003_sig0000006f,
      I2 => blk00000003_sig00000033,
      O => blk00000003_sig0000010e
    );
  blk00000003_blk00000147 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000000e6,
      I1 => blk00000003_sig0000003a,
      O => blk00000003_sig000000c8
    );
  blk00000003_blk00000146 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000000df,
      I1 => blk00000003_sig00000070,
      I2 => blk00000003_sig0000003a,
      O => blk00000003_sig000000cb
    );
  blk00000003_blk00000145 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000000e0,
      I1 => blk00000003_sig00000071,
      I2 => blk00000003_sig0000003a,
      O => blk00000003_sig000000ce
    );
  blk00000003_blk00000144 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000000e1,
      I1 => blk00000003_sig00000072,
      I2 => blk00000003_sig0000003a,
      O => blk00000003_sig000000d1
    );
  blk00000003_blk00000143 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000000e2,
      I1 => blk00000003_sig00000073,
      I2 => blk00000003_sig0000003a,
      O => blk00000003_sig000000d4
    );
  blk00000003_blk00000142 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000000e3,
      I1 => blk00000003_sig00000074,
      I2 => blk00000003_sig0000003a,
      O => blk00000003_sig000000d7
    );
  blk00000003_blk00000141 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000000e4,
      I1 => blk00000003_sig00000075,
      I2 => blk00000003_sig0000003a,
      O => blk00000003_sig000000da
    );
  blk00000003_blk00000140 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000000e5,
      I1 => blk00000003_sig00000076,
      I2 => blk00000003_sig0000003a,
      O => blk00000003_sig000000dd
    );
  blk00000003_blk0000013f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000040,
      I1 => blk00000003_sig00000077,
      I2 => blk00000003_sig0000003a,
      O => blk00000003_sig000000e9
    );
  blk00000003_blk0000013e : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000000c1,
      I1 => blk00000003_sig00000041,
      O => blk00000003_sig000000a3
    );
  blk00000003_blk0000013d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000000ba,
      I1 => blk00000003_sig00000078,
      I2 => blk00000003_sig00000041,
      O => blk00000003_sig000000a6
    );
  blk00000003_blk0000013c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000000bb,
      I1 => blk00000003_sig00000079,
      I2 => blk00000003_sig00000041,
      O => blk00000003_sig000000a9
    );
  blk00000003_blk0000013b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000000bc,
      I1 => blk00000003_sig0000007a,
      I2 => blk00000003_sig00000041,
      O => blk00000003_sig000000ac
    );
  blk00000003_blk0000013a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000000bd,
      I1 => blk00000003_sig0000007b,
      I2 => blk00000003_sig00000041,
      O => blk00000003_sig000000af
    );
  blk00000003_blk00000139 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000000be,
      I1 => blk00000003_sig0000007c,
      I2 => blk00000003_sig00000041,
      O => blk00000003_sig000000b2
    );
  blk00000003_blk00000138 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000000bf,
      I1 => blk00000003_sig0000007d,
      I2 => blk00000003_sig00000041,
      O => blk00000003_sig000000b5
    );
  blk00000003_blk00000137 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000000c0,
      I1 => blk00000003_sig0000007e,
      I2 => blk00000003_sig00000041,
      O => blk00000003_sig000000b8
    );
  blk00000003_blk00000136 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000047,
      I1 => blk00000003_sig0000007f,
      I2 => blk00000003_sig00000041,
      O => blk00000003_sig000000c4
    );
  blk00000003_blk00000135 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000049,
      I1 => blk00000003_sig00000087,
      O => blk00000003_sig0000009f
    );
  blk00000003_blk00000134 : LUT1
    generic map(
      INIT => X"1"
    )
    port map (
      I0 => blk00000003_sig0000015b,
      O => blk00000003_sig0000004a
    );
  blk00000003_blk00000133 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000185,
      Q => fractional(0)
    );
  blk00000003_blk00000132 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000178,
      Q => fractional(1)
    );
  blk00000003_blk00000131 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000175,
      Q => fractional(2)
    );
  blk00000003_blk00000130 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000172,
      Q => fractional(3)
    );
  blk00000003_blk0000012f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000016f,
      Q => fractional(4)
    );
  blk00000003_blk0000012e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000016c,
      Q => fractional(5)
    );
  blk00000003_blk0000012d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000169,
      Q => fractional(6)
    );
  blk00000003_blk0000012c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000166,
      Q => fractional(7)
    );
  blk00000003_blk0000012b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000017a,
      Q => blk00000003_sig00000188
    );
  blk00000003_blk0000012a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000017c,
      Q => blk00000003_sig00000187
    );
  blk00000003_blk00000129 : MULT_AND
    port map (
      I0 => blk00000003_sig0000005f,
      I1 => blk00000003_sig0000015b,
      LO => blk00000003_sig00000186
    );
  blk00000003_blk00000128 : MULT_AND
    port map (
      I0 => blk00000003_sig0000005d,
      I1 => blk00000003_sig0000015b,
      LO => blk00000003_sig00000183
    );
  blk00000003_blk00000127 : MULT_AND
    port map (
      I0 => blk00000003_sig0000005b,
      I1 => blk00000003_sig0000015b,
      LO => blk00000003_sig00000182
    );
  blk00000003_blk00000126 : MULT_AND
    port map (
      I0 => blk00000003_sig00000059,
      I1 => blk00000003_sig0000015b,
      LO => blk00000003_sig00000181
    );
  blk00000003_blk00000125 : MULT_AND
    port map (
      I0 => blk00000003_sig00000057,
      I1 => blk00000003_sig0000015b,
      LO => blk00000003_sig00000180
    );
  blk00000003_blk00000124 : MULT_AND
    port map (
      I0 => blk00000003_sig00000055,
      I1 => blk00000003_sig0000015b,
      LO => blk00000003_sig0000017f
    );
  blk00000003_blk00000123 : MULT_AND
    port map (
      I0 => blk00000003_sig00000053,
      I1 => blk00000003_sig0000015b,
      LO => blk00000003_sig0000017e
    );
  blk00000003_blk00000122 : MULT_AND
    port map (
      I0 => blk00000003_sig00000051,
      I1 => blk00000003_sig0000015b,
      LO => blk00000003_sig0000017d
    );
  blk00000003_blk00000121 : MULT_AND
    port map (
      I0 => blk00000003_sig0000001f,
      I1 => blk00000003_sig0000015b,
      LO => blk00000003_sig0000017b
    );
  blk00000003_blk00000120 : MUXCY
    port map (
      CI => blk00000003_sig0000001f,
      DI => blk00000003_sig00000186,
      S => blk00000003_sig00000184,
      O => blk00000003_sig00000176
    );
  blk00000003_blk0000011f : XORCY
    port map (
      CI => blk00000003_sig0000001f,
      LI => blk00000003_sig00000184,
      O => blk00000003_sig00000185
    );
  blk00000003_blk0000011e : MUXCY
    port map (
      CI => blk00000003_sig00000176,
      DI => blk00000003_sig00000183,
      S => blk00000003_sig00000177,
      O => blk00000003_sig00000173
    );
  blk00000003_blk0000011d : MUXCY
    port map (
      CI => blk00000003_sig00000173,
      DI => blk00000003_sig00000182,
      S => blk00000003_sig00000174,
      O => blk00000003_sig00000170
    );
  blk00000003_blk0000011c : MUXCY
    port map (
      CI => blk00000003_sig00000170,
      DI => blk00000003_sig00000181,
      S => blk00000003_sig00000171,
      O => blk00000003_sig0000016d
    );
  blk00000003_blk0000011b : MUXCY
    port map (
      CI => blk00000003_sig0000016d,
      DI => blk00000003_sig00000180,
      S => blk00000003_sig0000016e,
      O => blk00000003_sig0000016a
    );
  blk00000003_blk0000011a : MUXCY
    port map (
      CI => blk00000003_sig0000016a,
      DI => blk00000003_sig0000017f,
      S => blk00000003_sig0000016b,
      O => blk00000003_sig00000167
    );
  blk00000003_blk00000119 : MUXCY
    port map (
      CI => blk00000003_sig00000167,
      DI => blk00000003_sig0000017e,
      S => blk00000003_sig00000168,
      O => blk00000003_sig00000164
    );
  blk00000003_blk00000118 : MUXCY
    port map (
      CI => blk00000003_sig00000164,
      DI => blk00000003_sig0000017d,
      S => blk00000003_sig00000165,
      O => blk00000003_sig00000179
    );
  blk00000003_blk00000117 : MUXCY
    port map (
      CI => blk00000003_sig00000179,
      DI => blk00000003_sig0000017b,
      S => blk00000003_sig0000001f,
      O => blk00000003_sig0000017c
    );
  blk00000003_blk00000116 : XORCY
    port map (
      CI => blk00000003_sig00000179,
      LI => blk00000003_sig0000001f,
      O => blk00000003_sig0000017a
    );
  blk00000003_blk00000115 : XORCY
    port map (
      CI => blk00000003_sig00000176,
      LI => blk00000003_sig00000177,
      O => blk00000003_sig00000178
    );
  blk00000003_blk00000114 : XORCY
    port map (
      CI => blk00000003_sig00000173,
      LI => blk00000003_sig00000174,
      O => blk00000003_sig00000175
    );
  blk00000003_blk00000113 : XORCY
    port map (
      CI => blk00000003_sig00000170,
      LI => blk00000003_sig00000171,
      O => blk00000003_sig00000172
    );
  blk00000003_blk00000112 : XORCY
    port map (
      CI => blk00000003_sig0000016d,
      LI => blk00000003_sig0000016e,
      O => blk00000003_sig0000016f
    );
  blk00000003_blk00000111 : XORCY
    port map (
      CI => blk00000003_sig0000016a,
      LI => blk00000003_sig0000016b,
      O => blk00000003_sig0000016c
    );
  blk00000003_blk00000110 : XORCY
    port map (
      CI => blk00000003_sig00000167,
      LI => blk00000003_sig00000168,
      O => blk00000003_sig00000169
    );
  blk00000003_blk0000010f : XORCY
    port map (
      CI => blk00000003_sig00000164,
      LI => blk00000003_sig00000165,
      O => blk00000003_sig00000166
    );
  blk00000003_blk0000010e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a0,
      Q => blk00000003_sig000000c0
    );
  blk00000003_blk0000010d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000009d,
      Q => blk00000003_sig000000bf
    );
  blk00000003_blk0000010c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000009a,
      Q => blk00000003_sig000000be
    );
  blk00000003_blk0000010b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000097,
      Q => blk00000003_sig000000bd
    );
  blk00000003_blk0000010a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000094,
      Q => blk00000003_sig000000bc
    );
  blk00000003_blk00000109 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000091,
      Q => blk00000003_sig000000bb
    );
  blk00000003_blk00000108 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000008e,
      Q => blk00000003_sig000000ba
    );
  blk00000003_blk00000107 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000008b,
      Q => blk00000003_sig000000c1
    );
  blk00000003_blk00000106 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c5,
      Q => blk00000003_sig000000e5
    );
  blk00000003_blk00000105 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b9,
      Q => blk00000003_sig000000e4
    );
  blk00000003_blk00000104 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b6,
      Q => blk00000003_sig000000e3
    );
  blk00000003_blk00000103 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b3,
      Q => blk00000003_sig000000e2
    );
  blk00000003_blk00000102 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b0,
      Q => blk00000003_sig000000e1
    );
  blk00000003_blk00000101 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ad,
      Q => blk00000003_sig000000e0
    );
  blk00000003_blk00000100 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000aa,
      Q => blk00000003_sig000000df
    );
  blk00000003_blk000000ff : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a7,
      Q => blk00000003_sig000000e6
    );
  blk00000003_blk000000fe : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a4,
      Q => blk00000003_sig0000003a
    );
  blk00000003_blk000000fd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ea,
      Q => blk00000003_sig0000010a
    );
  blk00000003_blk000000fc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000de,
      Q => blk00000003_sig00000109
    );
  blk00000003_blk000000fb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000db,
      Q => blk00000003_sig00000108
    );
  blk00000003_blk000000fa : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d8,
      Q => blk00000003_sig00000107
    );
  blk00000003_blk000000f9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d5,
      Q => blk00000003_sig00000106
    );
  blk00000003_blk000000f8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d2,
      Q => blk00000003_sig00000105
    );
  blk00000003_blk000000f7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000cf,
      Q => blk00000003_sig00000104
    );
  blk00000003_blk000000f6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000cc,
      Q => blk00000003_sig0000010b
    );
  blk00000003_blk000000f5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c9,
      Q => blk00000003_sig00000033
    );
  blk00000003_blk000000f4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000010f,
      Q => blk00000003_sig0000012f
    );
  blk00000003_blk000000f3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000103,
      Q => blk00000003_sig0000012e
    );
  blk00000003_blk000000f2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000100,
      Q => blk00000003_sig0000012d
    );
  blk00000003_blk000000f1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000fd,
      Q => blk00000003_sig0000012c
    );
  blk00000003_blk000000f0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000fa,
      Q => blk00000003_sig0000012b
    );
  blk00000003_blk000000ef : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f7,
      Q => blk00000003_sig0000012a
    );
  blk00000003_blk000000ee : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f4,
      Q => blk00000003_sig00000129
    );
  blk00000003_blk000000ed : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f1,
      Q => blk00000003_sig00000130
    );
  blk00000003_blk000000ec : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ee,
      Q => blk00000003_sig0000002b
    );
  blk00000003_blk000000eb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000134,
      Q => blk00000003_sig00000154
    );
  blk00000003_blk000000ea : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000128,
      Q => blk00000003_sig00000153
    );
  blk00000003_blk000000e9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000125,
      Q => blk00000003_sig00000152
    );
  blk00000003_blk000000e8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000122,
      Q => blk00000003_sig00000151
    );
  blk00000003_blk000000e7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000011f,
      Q => blk00000003_sig00000150
    );
  blk00000003_blk000000e6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000011c,
      Q => blk00000003_sig0000014f
    );
  blk00000003_blk000000e5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000119,
      Q => blk00000003_sig0000014e
    );
  blk00000003_blk000000e4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000116,
      Q => blk00000003_sig00000155
    );
  blk00000003_blk000000e3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000113,
      Q => blk00000003_sig00000021
    );
  blk00000003_blk000000e2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000159,
      Q => blk00000003_sig00000163
    );
  blk00000003_blk000000e1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000014d,
      Q => blk00000003_sig00000162
    );
  blk00000003_blk000000e0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000014a,
      Q => blk00000003_sig00000161
    );
  blk00000003_blk000000df : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000147,
      Q => blk00000003_sig00000160
    );
  blk00000003_blk000000de : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000144,
      Q => blk00000003_sig0000015f
    );
  blk00000003_blk000000dd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000141,
      Q => blk00000003_sig0000015e
    );
  blk00000003_blk000000dc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000013e,
      Q => blk00000003_sig0000015d
    );
  blk00000003_blk000000db : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000013b,
      Q => blk00000003_sig0000015c
    );
  blk00000003_blk000000da : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000138,
      Q => blk00000003_sig0000015b
    );
  blk00000003_blk000000d9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000156,
      Q => blk00000003_sig0000015a
    );
  blk00000003_blk000000d8 : MUXCY
    port map (
      CI => blk00000003_sig00000157,
      DI => blk00000003_sig00000048,
      S => blk00000003_sig00000158,
      O => blk00000003_sig0000014b
    );
  blk00000003_blk000000d7 : XORCY
    port map (
      CI => blk00000003_sig00000157,
      LI => blk00000003_sig00000158,
      O => blk00000003_sig00000159
    );
  blk00000003_blk000000d6 : MUXCY
    port map (
      CI => blk00000003_sig00000136,
      DI => blk00000003_sig00000155,
      S => blk00000003_sig00000137,
      O => blk00000003_sig00000156
    );
  blk00000003_blk000000d5 : MUXCY
    port map (
      CI => blk00000003_sig0000014b,
      DI => blk00000003_sig00000154,
      S => blk00000003_sig0000014c,
      O => blk00000003_sig00000148
    );
  blk00000003_blk000000d4 : MUXCY
    port map (
      CI => blk00000003_sig00000148,
      DI => blk00000003_sig00000153,
      S => blk00000003_sig00000149,
      O => blk00000003_sig00000145
    );
  blk00000003_blk000000d3 : MUXCY
    port map (
      CI => blk00000003_sig00000145,
      DI => blk00000003_sig00000152,
      S => blk00000003_sig00000146,
      O => blk00000003_sig00000142
    );
  blk00000003_blk000000d2 : MUXCY
    port map (
      CI => blk00000003_sig00000142,
      DI => blk00000003_sig00000151,
      S => blk00000003_sig00000143,
      O => blk00000003_sig0000013f
    );
  blk00000003_blk000000d1 : MUXCY
    port map (
      CI => blk00000003_sig0000013f,
      DI => blk00000003_sig00000150,
      S => blk00000003_sig00000140,
      O => blk00000003_sig0000013c
    );
  blk00000003_blk000000d0 : MUXCY
    port map (
      CI => blk00000003_sig0000013c,
      DI => blk00000003_sig0000014f,
      S => blk00000003_sig0000013d,
      O => blk00000003_sig00000139
    );
  blk00000003_blk000000cf : MUXCY
    port map (
      CI => blk00000003_sig00000139,
      DI => blk00000003_sig0000014e,
      S => blk00000003_sig0000013a,
      O => blk00000003_sig00000136
    );
  blk00000003_blk000000ce : XORCY
    port map (
      CI => blk00000003_sig0000014b,
      LI => blk00000003_sig0000014c,
      O => blk00000003_sig0000014d
    );
  blk00000003_blk000000cd : XORCY
    port map (
      CI => blk00000003_sig00000148,
      LI => blk00000003_sig00000149,
      O => blk00000003_sig0000014a
    );
  blk00000003_blk000000cc : XORCY
    port map (
      CI => blk00000003_sig00000145,
      LI => blk00000003_sig00000146,
      O => blk00000003_sig00000147
    );
  blk00000003_blk000000cb : XORCY
    port map (
      CI => blk00000003_sig00000142,
      LI => blk00000003_sig00000143,
      O => blk00000003_sig00000144
    );
  blk00000003_blk000000ca : XORCY
    port map (
      CI => blk00000003_sig0000013f,
      LI => blk00000003_sig00000140,
      O => blk00000003_sig00000141
    );
  blk00000003_blk000000c9 : XORCY
    port map (
      CI => blk00000003_sig0000013c,
      LI => blk00000003_sig0000013d,
      O => blk00000003_sig0000013e
    );
  blk00000003_blk000000c8 : XORCY
    port map (
      CI => blk00000003_sig00000139,
      LI => blk00000003_sig0000013a,
      O => blk00000003_sig0000013b
    );
  blk00000003_blk000000c7 : XORCY
    port map (
      CI => blk00000003_sig00000136,
      LI => blk00000003_sig00000137,
      O => blk00000003_sig00000138
    );
  blk00000003_blk000000c6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000131,
      Q => blk00000003_sig00000135
    );
  blk00000003_blk000000c5 : MUXCY
    port map (
      CI => blk00000003_sig00000132,
      DI => blk00000003_sig00000032,
      S => blk00000003_sig00000133,
      O => blk00000003_sig00000126
    );
  blk00000003_blk000000c4 : XORCY
    port map (
      CI => blk00000003_sig00000132,
      LI => blk00000003_sig00000133,
      O => blk00000003_sig00000134
    );
  blk00000003_blk000000c3 : MUXCY
    port map (
      CI => blk00000003_sig00000111,
      DI => blk00000003_sig00000130,
      S => blk00000003_sig00000112,
      O => blk00000003_sig00000131
    );
  blk00000003_blk000000c2 : MUXCY
    port map (
      CI => blk00000003_sig00000126,
      DI => blk00000003_sig0000012f,
      S => blk00000003_sig00000127,
      O => blk00000003_sig00000123
    );
  blk00000003_blk000000c1 : MUXCY
    port map (
      CI => blk00000003_sig00000123,
      DI => blk00000003_sig0000012e,
      S => blk00000003_sig00000124,
      O => blk00000003_sig00000120
    );
  blk00000003_blk000000c0 : MUXCY
    port map (
      CI => blk00000003_sig00000120,
      DI => blk00000003_sig0000012d,
      S => blk00000003_sig00000121,
      O => blk00000003_sig0000011d
    );
  blk00000003_blk000000bf : MUXCY
    port map (
      CI => blk00000003_sig0000011d,
      DI => blk00000003_sig0000012c,
      S => blk00000003_sig0000011e,
      O => blk00000003_sig0000011a
    );
  blk00000003_blk000000be : MUXCY
    port map (
      CI => blk00000003_sig0000011a,
      DI => blk00000003_sig0000012b,
      S => blk00000003_sig0000011b,
      O => blk00000003_sig00000117
    );
  blk00000003_blk000000bd : MUXCY
    port map (
      CI => blk00000003_sig00000117,
      DI => blk00000003_sig0000012a,
      S => blk00000003_sig00000118,
      O => blk00000003_sig00000114
    );
  blk00000003_blk000000bc : MUXCY
    port map (
      CI => blk00000003_sig00000114,
      DI => blk00000003_sig00000129,
      S => blk00000003_sig00000115,
      O => blk00000003_sig00000111
    );
  blk00000003_blk000000bb : XORCY
    port map (
      CI => blk00000003_sig00000126,
      LI => blk00000003_sig00000127,
      O => blk00000003_sig00000128
    );
  blk00000003_blk000000ba : XORCY
    port map (
      CI => blk00000003_sig00000123,
      LI => blk00000003_sig00000124,
      O => blk00000003_sig00000125
    );
  blk00000003_blk000000b9 : XORCY
    port map (
      CI => blk00000003_sig00000120,
      LI => blk00000003_sig00000121,
      O => blk00000003_sig00000122
    );
  blk00000003_blk000000b8 : XORCY
    port map (
      CI => blk00000003_sig0000011d,
      LI => blk00000003_sig0000011e,
      O => blk00000003_sig0000011f
    );
  blk00000003_blk000000b7 : XORCY
    port map (
      CI => blk00000003_sig0000011a,
      LI => blk00000003_sig0000011b,
      O => blk00000003_sig0000011c
    );
  blk00000003_blk000000b6 : XORCY
    port map (
      CI => blk00000003_sig00000117,
      LI => blk00000003_sig00000118,
      O => blk00000003_sig00000119
    );
  blk00000003_blk000000b5 : XORCY
    port map (
      CI => blk00000003_sig00000114,
      LI => blk00000003_sig00000115,
      O => blk00000003_sig00000116
    );
  blk00000003_blk000000b4 : XORCY
    port map (
      CI => blk00000003_sig00000111,
      LI => blk00000003_sig00000112,
      O => blk00000003_sig00000113
    );
  blk00000003_blk000000b3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000010c,
      Q => blk00000003_sig00000110
    );
  blk00000003_blk000000b2 : MUXCY
    port map (
      CI => blk00000003_sig0000010d,
      DI => blk00000003_sig00000039,
      S => blk00000003_sig0000010e,
      O => blk00000003_sig00000101
    );
  blk00000003_blk000000b1 : XORCY
    port map (
      CI => blk00000003_sig0000010d,
      LI => blk00000003_sig0000010e,
      O => blk00000003_sig0000010f
    );
  blk00000003_blk000000b0 : MUXCY
    port map (
      CI => blk00000003_sig000000ec,
      DI => blk00000003_sig0000010b,
      S => blk00000003_sig000000ed,
      O => blk00000003_sig0000010c
    );
  blk00000003_blk000000af : MUXCY
    port map (
      CI => blk00000003_sig00000101,
      DI => blk00000003_sig0000010a,
      S => blk00000003_sig00000102,
      O => blk00000003_sig000000fe
    );
  blk00000003_blk000000ae : MUXCY
    port map (
      CI => blk00000003_sig000000fe,
      DI => blk00000003_sig00000109,
      S => blk00000003_sig000000ff,
      O => blk00000003_sig000000fb
    );
  blk00000003_blk000000ad : MUXCY
    port map (
      CI => blk00000003_sig000000fb,
      DI => blk00000003_sig00000108,
      S => blk00000003_sig000000fc,
      O => blk00000003_sig000000f8
    );
  blk00000003_blk000000ac : MUXCY
    port map (
      CI => blk00000003_sig000000f8,
      DI => blk00000003_sig00000107,
      S => blk00000003_sig000000f9,
      O => blk00000003_sig000000f5
    );
  blk00000003_blk000000ab : MUXCY
    port map (
      CI => blk00000003_sig000000f5,
      DI => blk00000003_sig00000106,
      S => blk00000003_sig000000f6,
      O => blk00000003_sig000000f2
    );
  blk00000003_blk000000aa : MUXCY
    port map (
      CI => blk00000003_sig000000f2,
      DI => blk00000003_sig00000105,
      S => blk00000003_sig000000f3,
      O => blk00000003_sig000000ef
    );
  blk00000003_blk000000a9 : MUXCY
    port map (
      CI => blk00000003_sig000000ef,
      DI => blk00000003_sig00000104,
      S => blk00000003_sig000000f0,
      O => blk00000003_sig000000ec
    );
  blk00000003_blk000000a8 : XORCY
    port map (
      CI => blk00000003_sig00000101,
      LI => blk00000003_sig00000102,
      O => blk00000003_sig00000103
    );
  blk00000003_blk000000a7 : XORCY
    port map (
      CI => blk00000003_sig000000fe,
      LI => blk00000003_sig000000ff,
      O => blk00000003_sig00000100
    );
  blk00000003_blk000000a6 : XORCY
    port map (
      CI => blk00000003_sig000000fb,
      LI => blk00000003_sig000000fc,
      O => blk00000003_sig000000fd
    );
  blk00000003_blk000000a5 : XORCY
    port map (
      CI => blk00000003_sig000000f8,
      LI => blk00000003_sig000000f9,
      O => blk00000003_sig000000fa
    );
  blk00000003_blk000000a4 : XORCY
    port map (
      CI => blk00000003_sig000000f5,
      LI => blk00000003_sig000000f6,
      O => blk00000003_sig000000f7
    );
  blk00000003_blk000000a3 : XORCY
    port map (
      CI => blk00000003_sig000000f2,
      LI => blk00000003_sig000000f3,
      O => blk00000003_sig000000f4
    );
  blk00000003_blk000000a2 : XORCY
    port map (
      CI => blk00000003_sig000000ef,
      LI => blk00000003_sig000000f0,
      O => blk00000003_sig000000f1
    );
  blk00000003_blk000000a1 : XORCY
    port map (
      CI => blk00000003_sig000000ec,
      LI => blk00000003_sig000000ed,
      O => blk00000003_sig000000ee
    );
  blk00000003_blk000000a0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e7,
      Q => blk00000003_sig000000eb
    );
  blk00000003_blk0000009f : MUXCY
    port map (
      CI => blk00000003_sig000000e8,
      DI => blk00000003_sig00000040,
      S => blk00000003_sig000000e9,
      O => blk00000003_sig000000dc
    );
  blk00000003_blk0000009e : XORCY
    port map (
      CI => blk00000003_sig000000e8,
      LI => blk00000003_sig000000e9,
      O => blk00000003_sig000000ea
    );
  blk00000003_blk0000009d : MUXCY
    port map (
      CI => blk00000003_sig000000c7,
      DI => blk00000003_sig000000e6,
      S => blk00000003_sig000000c8,
      O => blk00000003_sig000000e7
    );
  blk00000003_blk0000009c : MUXCY
    port map (
      CI => blk00000003_sig000000dc,
      DI => blk00000003_sig000000e5,
      S => blk00000003_sig000000dd,
      O => blk00000003_sig000000d9
    );
  blk00000003_blk0000009b : MUXCY
    port map (
      CI => blk00000003_sig000000d9,
      DI => blk00000003_sig000000e4,
      S => blk00000003_sig000000da,
      O => blk00000003_sig000000d6
    );
  blk00000003_blk0000009a : MUXCY
    port map (
      CI => blk00000003_sig000000d6,
      DI => blk00000003_sig000000e3,
      S => blk00000003_sig000000d7,
      O => blk00000003_sig000000d3
    );
  blk00000003_blk00000099 : MUXCY
    port map (
      CI => blk00000003_sig000000d3,
      DI => blk00000003_sig000000e2,
      S => blk00000003_sig000000d4,
      O => blk00000003_sig000000d0
    );
  blk00000003_blk00000098 : MUXCY
    port map (
      CI => blk00000003_sig000000d0,
      DI => blk00000003_sig000000e1,
      S => blk00000003_sig000000d1,
      O => blk00000003_sig000000cd
    );
  blk00000003_blk00000097 : MUXCY
    port map (
      CI => blk00000003_sig000000cd,
      DI => blk00000003_sig000000e0,
      S => blk00000003_sig000000ce,
      O => blk00000003_sig000000ca
    );
  blk00000003_blk00000096 : MUXCY
    port map (
      CI => blk00000003_sig000000ca,
      DI => blk00000003_sig000000df,
      S => blk00000003_sig000000cb,
      O => blk00000003_sig000000c7
    );
  blk00000003_blk00000095 : XORCY
    port map (
      CI => blk00000003_sig000000dc,
      LI => blk00000003_sig000000dd,
      O => blk00000003_sig000000de
    );
  blk00000003_blk00000094 : XORCY
    port map (
      CI => blk00000003_sig000000d9,
      LI => blk00000003_sig000000da,
      O => blk00000003_sig000000db
    );
  blk00000003_blk00000093 : XORCY
    port map (
      CI => blk00000003_sig000000d6,
      LI => blk00000003_sig000000d7,
      O => blk00000003_sig000000d8
    );
  blk00000003_blk00000092 : XORCY
    port map (
      CI => blk00000003_sig000000d3,
      LI => blk00000003_sig000000d4,
      O => blk00000003_sig000000d5
    );
  blk00000003_blk00000091 : XORCY
    port map (
      CI => blk00000003_sig000000d0,
      LI => blk00000003_sig000000d1,
      O => blk00000003_sig000000d2
    );
  blk00000003_blk00000090 : XORCY
    port map (
      CI => blk00000003_sig000000cd,
      LI => blk00000003_sig000000ce,
      O => blk00000003_sig000000cf
    );
  blk00000003_blk0000008f : XORCY
    port map (
      CI => blk00000003_sig000000ca,
      LI => blk00000003_sig000000cb,
      O => blk00000003_sig000000cc
    );
  blk00000003_blk0000008e : XORCY
    port map (
      CI => blk00000003_sig000000c7,
      LI => blk00000003_sig000000c8,
      O => blk00000003_sig000000c9
    );
  blk00000003_blk0000008d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c2,
      Q => blk00000003_sig000000c6
    );
  blk00000003_blk0000008c : MUXCY
    port map (
      CI => blk00000003_sig000000c3,
      DI => blk00000003_sig00000047,
      S => blk00000003_sig000000c4,
      O => blk00000003_sig000000b7
    );
  blk00000003_blk0000008b : XORCY
    port map (
      CI => blk00000003_sig000000c3,
      LI => blk00000003_sig000000c4,
      O => blk00000003_sig000000c5
    );
  blk00000003_blk0000008a : MUXCY
    port map (
      CI => blk00000003_sig000000a2,
      DI => blk00000003_sig000000c1,
      S => blk00000003_sig000000a3,
      O => blk00000003_sig000000c2
    );
  blk00000003_blk00000089 : MUXCY
    port map (
      CI => blk00000003_sig000000b7,
      DI => blk00000003_sig000000c0,
      S => blk00000003_sig000000b8,
      O => blk00000003_sig000000b4
    );
  blk00000003_blk00000088 : MUXCY
    port map (
      CI => blk00000003_sig000000b4,
      DI => blk00000003_sig000000bf,
      S => blk00000003_sig000000b5,
      O => blk00000003_sig000000b1
    );
  blk00000003_blk00000087 : MUXCY
    port map (
      CI => blk00000003_sig000000b1,
      DI => blk00000003_sig000000be,
      S => blk00000003_sig000000b2,
      O => blk00000003_sig000000ae
    );
  blk00000003_blk00000086 : MUXCY
    port map (
      CI => blk00000003_sig000000ae,
      DI => blk00000003_sig000000bd,
      S => blk00000003_sig000000af,
      O => blk00000003_sig000000ab
    );
  blk00000003_blk00000085 : MUXCY
    port map (
      CI => blk00000003_sig000000ab,
      DI => blk00000003_sig000000bc,
      S => blk00000003_sig000000ac,
      O => blk00000003_sig000000a8
    );
  blk00000003_blk00000084 : MUXCY
    port map (
      CI => blk00000003_sig000000a8,
      DI => blk00000003_sig000000bb,
      S => blk00000003_sig000000a9,
      O => blk00000003_sig000000a5
    );
  blk00000003_blk00000083 : MUXCY
    port map (
      CI => blk00000003_sig000000a5,
      DI => blk00000003_sig000000ba,
      S => blk00000003_sig000000a6,
      O => blk00000003_sig000000a2
    );
  blk00000003_blk00000082 : XORCY
    port map (
      CI => blk00000003_sig000000b7,
      LI => blk00000003_sig000000b8,
      O => blk00000003_sig000000b9
    );
  blk00000003_blk00000081 : XORCY
    port map (
      CI => blk00000003_sig000000b4,
      LI => blk00000003_sig000000b5,
      O => blk00000003_sig000000b6
    );
  blk00000003_blk00000080 : XORCY
    port map (
      CI => blk00000003_sig000000b1,
      LI => blk00000003_sig000000b2,
      O => blk00000003_sig000000b3
    );
  blk00000003_blk0000007f : XORCY
    port map (
      CI => blk00000003_sig000000ae,
      LI => blk00000003_sig000000af,
      O => blk00000003_sig000000b0
    );
  blk00000003_blk0000007e : XORCY
    port map (
      CI => blk00000003_sig000000ab,
      LI => blk00000003_sig000000ac,
      O => blk00000003_sig000000ad
    );
  blk00000003_blk0000007d : XORCY
    port map (
      CI => blk00000003_sig000000a8,
      LI => blk00000003_sig000000a9,
      O => blk00000003_sig000000aa
    );
  blk00000003_blk0000007c : XORCY
    port map (
      CI => blk00000003_sig000000a5,
      LI => blk00000003_sig000000a6,
      O => blk00000003_sig000000a7
    );
  blk00000003_blk0000007b : XORCY
    port map (
      CI => blk00000003_sig000000a2,
      LI => blk00000003_sig000000a3,
      O => blk00000003_sig000000a4
    );
  blk00000003_blk0000007a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000009e,
      Q => blk00000003_sig000000a1
    );
  blk00000003_blk00000079 : MUXCY
    port map (
      CI => NlwRenamedSig_OI_rfd,
      DI => blk00000003_sig00000049,
      S => blk00000003_sig0000009f,
      O => blk00000003_sig0000009b
    );
  blk00000003_blk00000078 : XORCY
    port map (
      CI => NlwRenamedSig_OI_rfd,
      LI => blk00000003_sig0000009f,
      O => blk00000003_sig000000a0
    );
  blk00000003_blk00000077 : MUXCY
    port map (
      CI => blk00000003_sig00000088,
      DI => blk00000003_sig0000001f,
      S => NlwRenamedSig_OI_rfd,
      O => blk00000003_sig0000009e
    );
  blk00000003_blk00000076 : MUXCY
    port map (
      CI => blk00000003_sig0000009b,
      DI => blk00000003_sig0000001f,
      S => blk00000003_sig0000009c,
      O => blk00000003_sig00000098
    );
  blk00000003_blk00000075 : MUXCY
    port map (
      CI => blk00000003_sig00000098,
      DI => blk00000003_sig0000001f,
      S => blk00000003_sig00000099,
      O => blk00000003_sig00000095
    );
  blk00000003_blk00000074 : MUXCY
    port map (
      CI => blk00000003_sig00000095,
      DI => blk00000003_sig0000001f,
      S => blk00000003_sig00000096,
      O => blk00000003_sig00000092
    );
  blk00000003_blk00000073 : MUXCY
    port map (
      CI => blk00000003_sig00000092,
      DI => blk00000003_sig0000001f,
      S => blk00000003_sig00000093,
      O => blk00000003_sig0000008f
    );
  blk00000003_blk00000072 : MUXCY
    port map (
      CI => blk00000003_sig0000008f,
      DI => blk00000003_sig0000001f,
      S => blk00000003_sig00000090,
      O => blk00000003_sig0000008c
    );
  blk00000003_blk00000071 : MUXCY
    port map (
      CI => blk00000003_sig0000008c,
      DI => blk00000003_sig0000001f,
      S => blk00000003_sig0000008d,
      O => blk00000003_sig00000089
    );
  blk00000003_blk00000070 : MUXCY
    port map (
      CI => blk00000003_sig00000089,
      DI => blk00000003_sig0000001f,
      S => blk00000003_sig0000008a,
      O => blk00000003_sig00000088
    );
  blk00000003_blk0000006f : XORCY
    port map (
      CI => blk00000003_sig0000009b,
      LI => blk00000003_sig0000009c,
      O => blk00000003_sig0000009d
    );
  blk00000003_blk0000006e : XORCY
    port map (
      CI => blk00000003_sig00000098,
      LI => blk00000003_sig00000099,
      O => blk00000003_sig0000009a
    );
  blk00000003_blk0000006d : XORCY
    port map (
      CI => blk00000003_sig00000095,
      LI => blk00000003_sig00000096,
      O => blk00000003_sig00000097
    );
  blk00000003_blk0000006c : XORCY
    port map (
      CI => blk00000003_sig00000092,
      LI => blk00000003_sig00000093,
      O => blk00000003_sig00000094
    );
  blk00000003_blk0000006b : XORCY
    port map (
      CI => blk00000003_sig0000008f,
      LI => blk00000003_sig00000090,
      O => blk00000003_sig00000091
    );
  blk00000003_blk0000006a : XORCY
    port map (
      CI => blk00000003_sig0000008c,
      LI => blk00000003_sig0000008d,
      O => blk00000003_sig0000008e
    );
  blk00000003_blk00000069 : XORCY
    port map (
      CI => blk00000003_sig00000089,
      LI => blk00000003_sig0000008a,
      O => blk00000003_sig0000008b
    );
  blk00000003_blk00000068 : XORCY
    port map (
      CI => blk00000003_sig00000088,
      LI => NlwRenamedSig_OI_rfd,
      O => NLW_blk00000003_blk00000068_O_UNCONNECTED
    );
  blk00000003_blk00000067 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(0),
      Q => blk00000003_sig00000087
    );
  blk00000003_blk00000066 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(1),
      Q => blk00000003_sig00000086
    );
  blk00000003_blk00000065 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(2),
      Q => blk00000003_sig00000085
    );
  blk00000003_blk00000064 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(3),
      Q => blk00000003_sig00000084
    );
  blk00000003_blk00000063 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(4),
      Q => blk00000003_sig00000083
    );
  blk00000003_blk00000062 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(5),
      Q => blk00000003_sig00000082
    );
  blk00000003_blk00000061 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(6),
      Q => blk00000003_sig00000081
    );
  blk00000003_blk00000060 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(7),
      Q => blk00000003_sig00000080
    );
  blk00000003_blk0000005f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000087,
      Q => blk00000003_sig0000007f
    );
  blk00000003_blk0000005e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000086,
      Q => blk00000003_sig0000007e
    );
  blk00000003_blk0000005d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000085,
      Q => blk00000003_sig0000007d
    );
  blk00000003_blk0000005c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000084,
      Q => blk00000003_sig0000007c
    );
  blk00000003_blk0000005b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000083,
      Q => blk00000003_sig0000007b
    );
  blk00000003_blk0000005a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000082,
      Q => blk00000003_sig0000007a
    );
  blk00000003_blk00000059 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000081,
      Q => blk00000003_sig00000079
    );
  blk00000003_blk00000058 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000080,
      Q => blk00000003_sig00000078
    );
  blk00000003_blk00000057 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007f,
      Q => blk00000003_sig00000077
    );
  blk00000003_blk00000056 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007e,
      Q => blk00000003_sig00000076
    );
  blk00000003_blk00000055 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007d,
      Q => blk00000003_sig00000075
    );
  blk00000003_blk00000054 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007c,
      Q => blk00000003_sig00000074
    );
  blk00000003_blk00000053 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007b,
      Q => blk00000003_sig00000073
    );
  blk00000003_blk00000052 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007a,
      Q => blk00000003_sig00000072
    );
  blk00000003_blk00000051 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000079,
      Q => blk00000003_sig00000071
    );
  blk00000003_blk00000050 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000078,
      Q => blk00000003_sig00000070
    );
  blk00000003_blk0000004f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000077,
      Q => blk00000003_sig0000006f
    );
  blk00000003_blk0000004e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000076,
      Q => blk00000003_sig0000006e
    );
  blk00000003_blk0000004d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000075,
      Q => blk00000003_sig0000006d
    );
  blk00000003_blk0000004c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000074,
      Q => blk00000003_sig0000006c
    );
  blk00000003_blk0000004b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000073,
      Q => blk00000003_sig0000006b
    );
  blk00000003_blk0000004a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000072,
      Q => blk00000003_sig0000006a
    );
  blk00000003_blk00000049 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000071,
      Q => blk00000003_sig00000069
    );
  blk00000003_blk00000048 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000070,
      Q => blk00000003_sig00000068
    );
  blk00000003_blk00000047 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006f,
      Q => blk00000003_sig00000067
    );
  blk00000003_blk00000046 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006e,
      Q => blk00000003_sig00000066
    );
  blk00000003_blk00000045 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006d,
      Q => blk00000003_sig00000065
    );
  blk00000003_blk00000044 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006c,
      Q => blk00000003_sig00000064
    );
  blk00000003_blk00000043 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006b,
      Q => blk00000003_sig00000063
    );
  blk00000003_blk00000042 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006a,
      Q => blk00000003_sig00000062
    );
  blk00000003_blk00000041 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000069,
      Q => blk00000003_sig00000061
    );
  blk00000003_blk00000040 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000068,
      Q => blk00000003_sig00000060
    );
  blk00000003_blk0000003f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000067,
      Q => blk00000003_sig0000005e
    );
  blk00000003_blk0000003e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000066,
      Q => blk00000003_sig0000005c
    );
  blk00000003_blk0000003d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000065,
      Q => blk00000003_sig0000005a
    );
  blk00000003_blk0000003c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000064,
      Q => blk00000003_sig00000058
    );
  blk00000003_blk0000003b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000063,
      Q => blk00000003_sig00000056
    );
  blk00000003_blk0000003a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000062,
      Q => blk00000003_sig00000054
    );
  blk00000003_blk00000039 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000061,
      Q => blk00000003_sig00000052
    );
  blk00000003_blk00000038 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000060,
      Q => blk00000003_sig00000050
    );
  blk00000003_blk00000037 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000005e,
      Q => blk00000003_sig0000005f
    );
  blk00000003_blk00000036 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000005c,
      Q => blk00000003_sig0000005d
    );
  blk00000003_blk00000035 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000005a,
      Q => blk00000003_sig0000005b
    );
  blk00000003_blk00000034 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000058,
      Q => blk00000003_sig00000059
    );
  blk00000003_blk00000033 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000056,
      Q => blk00000003_sig00000057
    );
  blk00000003_blk00000032 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000054,
      Q => blk00000003_sig00000055
    );
  blk00000003_blk00000031 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000052,
      Q => blk00000003_sig00000053
    );
  blk00000003_blk00000030 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000050,
      Q => blk00000003_sig00000051
    );
  blk00000003_blk0000002f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000004f,
      Q => quotient(5)
    );
  blk00000003_blk0000002e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000004e,
      Q => quotient(4)
    );
  blk00000003_blk0000002d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000004d,
      Q => quotient(3)
    );
  blk00000003_blk0000002c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000004c,
      Q => quotient(2)
    );
  blk00000003_blk0000002b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000004b,
      Q => quotient(1)
    );
  blk00000003_blk0000002a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000004a,
      Q => quotient(0)
    );
  blk00000003_blk00000029 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(5),
      Q => blk00000003_sig00000049
    );
  blk00000003_blk00000028 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(4),
      Q => blk00000003_sig00000046
    );
  blk00000003_blk00000027 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(3),
      Q => blk00000003_sig00000045
    );
  blk00000003_blk00000026 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(2),
      Q => blk00000003_sig00000044
    );
  blk00000003_blk00000025 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(1),
      Q => blk00000003_sig00000043
    );
  blk00000003_blk00000024 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(0),
      Q => blk00000003_sig00000042
    );
  blk00000003_blk00000023 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000030,
      Q => blk00000003_sig00000048
    );
  blk00000003_blk00000022 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000046,
      Q => blk00000003_sig00000047
    );
  blk00000003_blk00000021 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000045,
      Q => blk00000003_sig0000003f
    );
  blk00000003_blk00000020 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000044,
      Q => blk00000003_sig0000003e
    );
  blk00000003_blk0000001f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000043,
      Q => blk00000003_sig0000003d
    );
  blk00000003_blk0000001e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000042,
      Q => blk00000003_sig0000003c
    );
  blk00000003_blk0000001d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000041,
      Q => blk00000003_sig0000003b
    );
  blk00000003_blk0000001c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000003f,
      Q => blk00000003_sig00000040
    );
  blk00000003_blk0000001b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000003e,
      Q => blk00000003_sig00000038
    );
  blk00000003_blk0000001a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000003d,
      Q => blk00000003_sig00000037
    );
  blk00000003_blk00000019 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000003c,
      Q => blk00000003_sig00000036
    );
  blk00000003_blk00000018 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000003b,
      Q => blk00000003_sig00000035
    );
  blk00000003_blk00000017 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000003a,
      Q => blk00000003_sig00000034
    );
  blk00000003_blk00000016 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000038,
      Q => blk00000003_sig00000039
    );
  blk00000003_blk00000015 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000037,
      Q => blk00000003_sig00000031
    );
  blk00000003_blk00000014 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000036,
      Q => blk00000003_sig0000002f
    );
  blk00000003_blk00000013 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000035,
      Q => blk00000003_sig0000002e
    );
  blk00000003_blk00000012 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000034,
      Q => blk00000003_sig0000002d
    );
  blk00000003_blk00000011 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000033,
      Q => blk00000003_sig0000002c
    );
  blk00000003_blk00000010 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000031,
      Q => blk00000003_sig00000032
    );
  blk00000003_blk0000000f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000002f,
      Q => blk00000003_sig00000030
    );
  blk00000003_blk0000000e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000002e,
      Q => blk00000003_sig00000029
    );
  blk00000003_blk0000000d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000002d,
      Q => blk00000003_sig00000027
    );
  blk00000003_blk0000000c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000002c,
      Q => blk00000003_sig00000025
    );
  blk00000003_blk0000000b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000002b,
      Q => blk00000003_sig00000023
    );
  blk00000003_blk0000000a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000029,
      Q => blk00000003_sig0000002a
    );
  blk00000003_blk00000009 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000027,
      Q => blk00000003_sig00000028
    );
  blk00000003_blk00000008 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000025,
      Q => blk00000003_sig00000026
    );
  blk00000003_blk00000007 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000023,
      Q => blk00000003_sig00000024
    );
  blk00000003_blk00000006 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000021,
      Q => blk00000003_sig00000022
    );
  blk00000003_blk00000005 : VCC
    port map (
      P => NlwRenamedSig_OI_rfd
    );
  blk00000003_blk00000004 : GND
    port map (
      G => blk00000003_sig0000001f
    );

end STRUCTURE;

-- synthesis translate_on
--------------------------------------------------------------------------------
-- Copyright (c) 1995-2011 Xilinx, Inc.  All rights reserved.
--------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version: O.61xd
--  \   \         Application: netgen
--  /   /         Filename: dv_gn_v3_0_56e83f20db65428d.vhd
-- /___/   /\     Timestamp: Mon Jul 23 19:55:53 2012
-- \   \  /  \ 
--  \___\/\___\
--             
-- Command	: -intstyle ise -w -sim -ofmt vhdl ./tmp/_cg/dv_gn_v3_0_56e83f20db65428d.ngc ./tmp/_cg/dv_gn_v3_0_56e83f20db65428d.vhd 
-- Device	: 6vcx75tff484-2
-- Input file	: ./tmp/_cg/dv_gn_v3_0_56e83f20db65428d.ngc
-- Output file	: ./tmp/_cg/dv_gn_v3_0_56e83f20db65428d.vhd
-- # of Entities	: 1
-- Design Name	: dv_gn_v3_0_56e83f20db65428d
-- Xilinx	: c:\xilinx\13.2\ise_ds\ise\
--             
-- Purpose:    
--     This VHDL netlist is a verification model and uses simulation 
--     primitives which may not represent the true implementation of the 
--     device, however the netlist is functionally correct and should not 
--     be modified. This file cannot be synthesized and should only be used 
--     with supported simulation tools.
--             
-- Reference:  
--     Command Line Tools User Guide, Chapter 23
--     Synthesis and Simulation Design Guide, Chapter 6
--             
--------------------------------------------------------------------------------


-- synthesis translate_off
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;
use UNISIM.VPKG.ALL;

entity dv_gn_v3_0_56e83f20db65428d is
  port (
    ce : in STD_LOGIC := 'X'; 
    rfd : out STD_LOGIC; 
    clk : in STD_LOGIC := 'X'; 
    dividend : in STD_LOGIC_VECTOR ( 31 downto 0 ); 
    quotient : out STD_LOGIC_VECTOR ( 31 downto 0 ); 
    divisor : in STD_LOGIC_VECTOR ( 7 downto 0 ); 
    fractional : out STD_LOGIC_VECTOR ( 7 downto 0 ) 
  );
end dv_gn_v3_0_56e83f20db65428d;

architecture STRUCTURE of dv_gn_v3_0_56e83f20db65428d is
  signal NlwRenamedSig_OI_rfd : STD_LOGIC; 
  signal blk00000003_sig00000a5e : STD_LOGIC; 
  signal blk00000003_sig00000a5d : STD_LOGIC; 
  signal blk00000003_sig00000a5c : STD_LOGIC; 
  signal blk00000003_sig00000a5b : STD_LOGIC; 
  signal blk00000003_sig00000a5a : STD_LOGIC; 
  signal blk00000003_sig00000a59 : STD_LOGIC; 
  signal blk00000003_sig00000a58 : STD_LOGIC; 
  signal blk00000003_sig00000a57 : STD_LOGIC; 
  signal blk00000003_sig00000a56 : STD_LOGIC; 
  signal blk00000003_sig00000a55 : STD_LOGIC; 
  signal blk00000003_sig00000a54 : STD_LOGIC; 
  signal blk00000003_sig00000a53 : STD_LOGIC; 
  signal blk00000003_sig00000a52 : STD_LOGIC; 
  signal blk00000003_sig00000a51 : STD_LOGIC; 
  signal blk00000003_sig00000a50 : STD_LOGIC; 
  signal blk00000003_sig00000a4f : STD_LOGIC; 
  signal blk00000003_sig00000a4e : STD_LOGIC; 
  signal blk00000003_sig00000a4d : STD_LOGIC; 
  signal blk00000003_sig00000a4c : STD_LOGIC; 
  signal blk00000003_sig00000a4b : STD_LOGIC; 
  signal blk00000003_sig00000a4a : STD_LOGIC; 
  signal blk00000003_sig00000a49 : STD_LOGIC; 
  signal blk00000003_sig00000a48 : STD_LOGIC; 
  signal blk00000003_sig00000a47 : STD_LOGIC; 
  signal blk00000003_sig00000a46 : STD_LOGIC; 
  signal blk00000003_sig00000a45 : STD_LOGIC; 
  signal blk00000003_sig00000a44 : STD_LOGIC; 
  signal blk00000003_sig00000a43 : STD_LOGIC; 
  signal blk00000003_sig00000a42 : STD_LOGIC; 
  signal blk00000003_sig00000a41 : STD_LOGIC; 
  signal blk00000003_sig00000a40 : STD_LOGIC; 
  signal blk00000003_sig00000a3f : STD_LOGIC; 
  signal blk00000003_sig00000a3e : STD_LOGIC; 
  signal blk00000003_sig00000a3d : STD_LOGIC; 
  signal blk00000003_sig00000a3c : STD_LOGIC; 
  signal blk00000003_sig00000a3b : STD_LOGIC; 
  signal blk00000003_sig00000a3a : STD_LOGIC; 
  signal blk00000003_sig00000a39 : STD_LOGIC; 
  signal blk00000003_sig00000a38 : STD_LOGIC; 
  signal blk00000003_sig00000a37 : STD_LOGIC; 
  signal blk00000003_sig00000a36 : STD_LOGIC; 
  signal blk00000003_sig00000a35 : STD_LOGIC; 
  signal blk00000003_sig00000a34 : STD_LOGIC; 
  signal blk00000003_sig00000a33 : STD_LOGIC; 
  signal blk00000003_sig00000a32 : STD_LOGIC; 
  signal blk00000003_sig00000a31 : STD_LOGIC; 
  signal blk00000003_sig00000a30 : STD_LOGIC; 
  signal blk00000003_sig00000a2f : STD_LOGIC; 
  signal blk00000003_sig00000a2e : STD_LOGIC; 
  signal blk00000003_sig00000a2d : STD_LOGIC; 
  signal blk00000003_sig00000a2c : STD_LOGIC; 
  signal blk00000003_sig00000a2b : STD_LOGIC; 
  signal blk00000003_sig00000a2a : STD_LOGIC; 
  signal blk00000003_sig00000a29 : STD_LOGIC; 
  signal blk00000003_sig00000a28 : STD_LOGIC; 
  signal blk00000003_sig00000a27 : STD_LOGIC; 
  signal blk00000003_sig00000a26 : STD_LOGIC; 
  signal blk00000003_sig00000a25 : STD_LOGIC; 
  signal blk00000003_sig00000a24 : STD_LOGIC; 
  signal blk00000003_sig00000a23 : STD_LOGIC; 
  signal blk00000003_sig00000a22 : STD_LOGIC; 
  signal blk00000003_sig00000a21 : STD_LOGIC; 
  signal blk00000003_sig00000a20 : STD_LOGIC; 
  signal blk00000003_sig00000a1f : STD_LOGIC; 
  signal blk00000003_sig00000a1e : STD_LOGIC; 
  signal blk00000003_sig00000a1d : STD_LOGIC; 
  signal blk00000003_sig00000a1c : STD_LOGIC; 
  signal blk00000003_sig00000a1b : STD_LOGIC; 
  signal blk00000003_sig00000a1a : STD_LOGIC; 
  signal blk00000003_sig00000a19 : STD_LOGIC; 
  signal blk00000003_sig00000a18 : STD_LOGIC; 
  signal blk00000003_sig00000a17 : STD_LOGIC; 
  signal blk00000003_sig00000a16 : STD_LOGIC; 
  signal blk00000003_sig00000a15 : STD_LOGIC; 
  signal blk00000003_sig00000a14 : STD_LOGIC; 
  signal blk00000003_sig00000a13 : STD_LOGIC; 
  signal blk00000003_sig00000a12 : STD_LOGIC; 
  signal blk00000003_sig00000a11 : STD_LOGIC; 
  signal blk00000003_sig00000a10 : STD_LOGIC; 
  signal blk00000003_sig00000a0f : STD_LOGIC; 
  signal blk00000003_sig00000a0e : STD_LOGIC; 
  signal blk00000003_sig00000a0d : STD_LOGIC; 
  signal blk00000003_sig00000a0c : STD_LOGIC; 
  signal blk00000003_sig00000a0b : STD_LOGIC; 
  signal blk00000003_sig00000a0a : STD_LOGIC; 
  signal blk00000003_sig00000a09 : STD_LOGIC; 
  signal blk00000003_sig00000a08 : STD_LOGIC; 
  signal blk00000003_sig00000a07 : STD_LOGIC; 
  signal blk00000003_sig00000a06 : STD_LOGIC; 
  signal blk00000003_sig00000a05 : STD_LOGIC; 
  signal blk00000003_sig00000a04 : STD_LOGIC; 
  signal blk00000003_sig00000a03 : STD_LOGIC; 
  signal blk00000003_sig00000a02 : STD_LOGIC; 
  signal blk00000003_sig00000a01 : STD_LOGIC; 
  signal blk00000003_sig00000a00 : STD_LOGIC; 
  signal blk00000003_sig000009ff : STD_LOGIC; 
  signal blk00000003_sig000009fe : STD_LOGIC; 
  signal blk00000003_sig000009fd : STD_LOGIC; 
  signal blk00000003_sig000009fc : STD_LOGIC; 
  signal blk00000003_sig000009fb : STD_LOGIC; 
  signal blk00000003_sig000009fa : STD_LOGIC; 
  signal blk00000003_sig000009f9 : STD_LOGIC; 
  signal blk00000003_sig000009f8 : STD_LOGIC; 
  signal blk00000003_sig000009f7 : STD_LOGIC; 
  signal blk00000003_sig000009f6 : STD_LOGIC; 
  signal blk00000003_sig000009f5 : STD_LOGIC; 
  signal blk00000003_sig000009f4 : STD_LOGIC; 
  signal blk00000003_sig000009f3 : STD_LOGIC; 
  signal blk00000003_sig000009f2 : STD_LOGIC; 
  signal blk00000003_sig000009f1 : STD_LOGIC; 
  signal blk00000003_sig000009f0 : STD_LOGIC; 
  signal blk00000003_sig000009ef : STD_LOGIC; 
  signal blk00000003_sig000009ee : STD_LOGIC; 
  signal blk00000003_sig000009ed : STD_LOGIC; 
  signal blk00000003_sig000009ec : STD_LOGIC; 
  signal blk00000003_sig000009eb : STD_LOGIC; 
  signal blk00000003_sig000009ea : STD_LOGIC; 
  signal blk00000003_sig000009e9 : STD_LOGIC; 
  signal blk00000003_sig000009e8 : STD_LOGIC; 
  signal blk00000003_sig000009e7 : STD_LOGIC; 
  signal blk00000003_sig000009e6 : STD_LOGIC; 
  signal blk00000003_sig000009e5 : STD_LOGIC; 
  signal blk00000003_sig000009e4 : STD_LOGIC; 
  signal blk00000003_sig000009e3 : STD_LOGIC; 
  signal blk00000003_sig000009e2 : STD_LOGIC; 
  signal blk00000003_sig000009e1 : STD_LOGIC; 
  signal blk00000003_sig000009e0 : STD_LOGIC; 
  signal blk00000003_sig000009df : STD_LOGIC; 
  signal blk00000003_sig000009de : STD_LOGIC; 
  signal blk00000003_sig000009dd : STD_LOGIC; 
  signal blk00000003_sig000009dc : STD_LOGIC; 
  signal blk00000003_sig000009db : STD_LOGIC; 
  signal blk00000003_sig000009da : STD_LOGIC; 
  signal blk00000003_sig000009d9 : STD_LOGIC; 
  signal blk00000003_sig000009d8 : STD_LOGIC; 
  signal blk00000003_sig000009d7 : STD_LOGIC; 
  signal blk00000003_sig000009d6 : STD_LOGIC; 
  signal blk00000003_sig000009d5 : STD_LOGIC; 
  signal blk00000003_sig000009d4 : STD_LOGIC; 
  signal blk00000003_sig000009d3 : STD_LOGIC; 
  signal blk00000003_sig000009d2 : STD_LOGIC; 
  signal blk00000003_sig000009d1 : STD_LOGIC; 
  signal blk00000003_sig000009d0 : STD_LOGIC; 
  signal blk00000003_sig000009cf : STD_LOGIC; 
  signal blk00000003_sig000009ce : STD_LOGIC; 
  signal blk00000003_sig000009cd : STD_LOGIC; 
  signal blk00000003_sig000009cc : STD_LOGIC; 
  signal blk00000003_sig000009cb : STD_LOGIC; 
  signal blk00000003_sig000009ca : STD_LOGIC; 
  signal blk00000003_sig000009c9 : STD_LOGIC; 
  signal blk00000003_sig000009c8 : STD_LOGIC; 
  signal blk00000003_sig000009c7 : STD_LOGIC; 
  signal blk00000003_sig000009c6 : STD_LOGIC; 
  signal blk00000003_sig000009c5 : STD_LOGIC; 
  signal blk00000003_sig000009c4 : STD_LOGIC; 
  signal blk00000003_sig000009c3 : STD_LOGIC; 
  signal blk00000003_sig000009c2 : STD_LOGIC; 
  signal blk00000003_sig000009c1 : STD_LOGIC; 
  signal blk00000003_sig000009c0 : STD_LOGIC; 
  signal blk00000003_sig000009bf : STD_LOGIC; 
  signal blk00000003_sig000009be : STD_LOGIC; 
  signal blk00000003_sig000009bd : STD_LOGIC; 
  signal blk00000003_sig000009bc : STD_LOGIC; 
  signal blk00000003_sig000009bb : STD_LOGIC; 
  signal blk00000003_sig000009ba : STD_LOGIC; 
  signal blk00000003_sig000009b9 : STD_LOGIC; 
  signal blk00000003_sig000009b8 : STD_LOGIC; 
  signal blk00000003_sig000009b7 : STD_LOGIC; 
  signal blk00000003_sig000009b6 : STD_LOGIC; 
  signal blk00000003_sig000009b5 : STD_LOGIC; 
  signal blk00000003_sig000009b4 : STD_LOGIC; 
  signal blk00000003_sig000009b3 : STD_LOGIC; 
  signal blk00000003_sig000009b2 : STD_LOGIC; 
  signal blk00000003_sig000009b1 : STD_LOGIC; 
  signal blk00000003_sig000009b0 : STD_LOGIC; 
  signal blk00000003_sig000009af : STD_LOGIC; 
  signal blk00000003_sig000009ae : STD_LOGIC; 
  signal blk00000003_sig000009ad : STD_LOGIC; 
  signal blk00000003_sig000009ac : STD_LOGIC; 
  signal blk00000003_sig000009ab : STD_LOGIC; 
  signal blk00000003_sig000009aa : STD_LOGIC; 
  signal blk00000003_sig000009a9 : STD_LOGIC; 
  signal blk00000003_sig000009a8 : STD_LOGIC; 
  signal blk00000003_sig000009a7 : STD_LOGIC; 
  signal blk00000003_sig000009a6 : STD_LOGIC; 
  signal blk00000003_sig000009a5 : STD_LOGIC; 
  signal blk00000003_sig000009a4 : STD_LOGIC; 
  signal blk00000003_sig000009a3 : STD_LOGIC; 
  signal blk00000003_sig000009a2 : STD_LOGIC; 
  signal blk00000003_sig000009a1 : STD_LOGIC; 
  signal blk00000003_sig000009a0 : STD_LOGIC; 
  signal blk00000003_sig0000099f : STD_LOGIC; 
  signal blk00000003_sig0000099e : STD_LOGIC; 
  signal blk00000003_sig0000099d : STD_LOGIC; 
  signal blk00000003_sig0000099c : STD_LOGIC; 
  signal blk00000003_sig0000099b : STD_LOGIC; 
  signal blk00000003_sig0000099a : STD_LOGIC; 
  signal blk00000003_sig00000999 : STD_LOGIC; 
  signal blk00000003_sig00000998 : STD_LOGIC; 
  signal blk00000003_sig00000997 : STD_LOGIC; 
  signal blk00000003_sig00000996 : STD_LOGIC; 
  signal blk00000003_sig00000995 : STD_LOGIC; 
  signal blk00000003_sig00000994 : STD_LOGIC; 
  signal blk00000003_sig00000993 : STD_LOGIC; 
  signal blk00000003_sig00000992 : STD_LOGIC; 
  signal blk00000003_sig00000991 : STD_LOGIC; 
  signal blk00000003_sig00000990 : STD_LOGIC; 
  signal blk00000003_sig0000098f : STD_LOGIC; 
  signal blk00000003_sig0000098e : STD_LOGIC; 
  signal blk00000003_sig0000098d : STD_LOGIC; 
  signal blk00000003_sig0000098c : STD_LOGIC; 
  signal blk00000003_sig0000098b : STD_LOGIC; 
  signal blk00000003_sig0000098a : STD_LOGIC; 
  signal blk00000003_sig00000989 : STD_LOGIC; 
  signal blk00000003_sig00000988 : STD_LOGIC; 
  signal blk00000003_sig00000987 : STD_LOGIC; 
  signal blk00000003_sig00000986 : STD_LOGIC; 
  signal blk00000003_sig00000985 : STD_LOGIC; 
  signal blk00000003_sig00000984 : STD_LOGIC; 
  signal blk00000003_sig00000983 : STD_LOGIC; 
  signal blk00000003_sig00000982 : STD_LOGIC; 
  signal blk00000003_sig00000981 : STD_LOGIC; 
  signal blk00000003_sig00000980 : STD_LOGIC; 
  signal blk00000003_sig0000097f : STD_LOGIC; 
  signal blk00000003_sig0000097e : STD_LOGIC; 
  signal blk00000003_sig0000097d : STD_LOGIC; 
  signal blk00000003_sig0000097c : STD_LOGIC; 
  signal blk00000003_sig0000097b : STD_LOGIC; 
  signal blk00000003_sig0000097a : STD_LOGIC; 
  signal blk00000003_sig00000979 : STD_LOGIC; 
  signal blk00000003_sig00000978 : STD_LOGIC; 
  signal blk00000003_sig00000977 : STD_LOGIC; 
  signal blk00000003_sig00000976 : STD_LOGIC; 
  signal blk00000003_sig00000975 : STD_LOGIC; 
  signal blk00000003_sig00000974 : STD_LOGIC; 
  signal blk00000003_sig00000973 : STD_LOGIC; 
  signal blk00000003_sig00000972 : STD_LOGIC; 
  signal blk00000003_sig00000971 : STD_LOGIC; 
  signal blk00000003_sig00000970 : STD_LOGIC; 
  signal blk00000003_sig0000096f : STD_LOGIC; 
  signal blk00000003_sig0000096e : STD_LOGIC; 
  signal blk00000003_sig0000096d : STD_LOGIC; 
  signal blk00000003_sig0000096c : STD_LOGIC; 
  signal blk00000003_sig0000096b : STD_LOGIC; 
  signal blk00000003_sig0000096a : STD_LOGIC; 
  signal blk00000003_sig00000969 : STD_LOGIC; 
  signal blk00000003_sig00000968 : STD_LOGIC; 
  signal blk00000003_sig00000967 : STD_LOGIC; 
  signal blk00000003_sig00000966 : STD_LOGIC; 
  signal blk00000003_sig00000965 : STD_LOGIC; 
  signal blk00000003_sig00000964 : STD_LOGIC; 
  signal blk00000003_sig00000963 : STD_LOGIC; 
  signal blk00000003_sig00000962 : STD_LOGIC; 
  signal blk00000003_sig00000961 : STD_LOGIC; 
  signal blk00000003_sig00000960 : STD_LOGIC; 
  signal blk00000003_sig0000095f : STD_LOGIC; 
  signal blk00000003_sig0000095e : STD_LOGIC; 
  signal blk00000003_sig0000095d : STD_LOGIC; 
  signal blk00000003_sig0000095c : STD_LOGIC; 
  signal blk00000003_sig0000095b : STD_LOGIC; 
  signal blk00000003_sig0000095a : STD_LOGIC; 
  signal blk00000003_sig00000959 : STD_LOGIC; 
  signal blk00000003_sig00000958 : STD_LOGIC; 
  signal blk00000003_sig00000957 : STD_LOGIC; 
  signal blk00000003_sig00000956 : STD_LOGIC; 
  signal blk00000003_sig00000955 : STD_LOGIC; 
  signal blk00000003_sig00000954 : STD_LOGIC; 
  signal blk00000003_sig00000953 : STD_LOGIC; 
  signal blk00000003_sig00000952 : STD_LOGIC; 
  signal blk00000003_sig00000951 : STD_LOGIC; 
  signal blk00000003_sig00000950 : STD_LOGIC; 
  signal blk00000003_sig0000094f : STD_LOGIC; 
  signal blk00000003_sig0000094e : STD_LOGIC; 
  signal blk00000003_sig0000094d : STD_LOGIC; 
  signal blk00000003_sig0000094c : STD_LOGIC; 
  signal blk00000003_sig0000094b : STD_LOGIC; 
  signal blk00000003_sig0000094a : STD_LOGIC; 
  signal blk00000003_sig00000949 : STD_LOGIC; 
  signal blk00000003_sig00000948 : STD_LOGIC; 
  signal blk00000003_sig00000947 : STD_LOGIC; 
  signal blk00000003_sig00000946 : STD_LOGIC; 
  signal blk00000003_sig00000945 : STD_LOGIC; 
  signal blk00000003_sig00000944 : STD_LOGIC; 
  signal blk00000003_sig00000943 : STD_LOGIC; 
  signal blk00000003_sig00000942 : STD_LOGIC; 
  signal blk00000003_sig00000941 : STD_LOGIC; 
  signal blk00000003_sig00000940 : STD_LOGIC; 
  signal blk00000003_sig0000093f : STD_LOGIC; 
  signal blk00000003_sig0000093e : STD_LOGIC; 
  signal blk00000003_sig0000093d : STD_LOGIC; 
  signal blk00000003_sig0000093c : STD_LOGIC; 
  signal blk00000003_sig0000093b : STD_LOGIC; 
  signal blk00000003_sig0000093a : STD_LOGIC; 
  signal blk00000003_sig00000939 : STD_LOGIC; 
  signal blk00000003_sig00000938 : STD_LOGIC; 
  signal blk00000003_sig00000937 : STD_LOGIC; 
  signal blk00000003_sig00000936 : STD_LOGIC; 
  signal blk00000003_sig00000935 : STD_LOGIC; 
  signal blk00000003_sig00000934 : STD_LOGIC; 
  signal blk00000003_sig00000933 : STD_LOGIC; 
  signal blk00000003_sig00000932 : STD_LOGIC; 
  signal blk00000003_sig00000931 : STD_LOGIC; 
  signal blk00000003_sig00000930 : STD_LOGIC; 
  signal blk00000003_sig0000092f : STD_LOGIC; 
  signal blk00000003_sig0000092e : STD_LOGIC; 
  signal blk00000003_sig0000092d : STD_LOGIC; 
  signal blk00000003_sig0000092c : STD_LOGIC; 
  signal blk00000003_sig0000092b : STD_LOGIC; 
  signal blk00000003_sig0000092a : STD_LOGIC; 
  signal blk00000003_sig00000929 : STD_LOGIC; 
  signal blk00000003_sig00000928 : STD_LOGIC; 
  signal blk00000003_sig00000927 : STD_LOGIC; 
  signal blk00000003_sig00000926 : STD_LOGIC; 
  signal blk00000003_sig00000925 : STD_LOGIC; 
  signal blk00000003_sig00000924 : STD_LOGIC; 
  signal blk00000003_sig00000923 : STD_LOGIC; 
  signal blk00000003_sig00000922 : STD_LOGIC; 
  signal blk00000003_sig00000921 : STD_LOGIC; 
  signal blk00000003_sig00000920 : STD_LOGIC; 
  signal blk00000003_sig0000091f : STD_LOGIC; 
  signal blk00000003_sig0000091e : STD_LOGIC; 
  signal blk00000003_sig0000091d : STD_LOGIC; 
  signal blk00000003_sig0000091c : STD_LOGIC; 
  signal blk00000003_sig0000091b : STD_LOGIC; 
  signal blk00000003_sig0000091a : STD_LOGIC; 
  signal blk00000003_sig00000919 : STD_LOGIC; 
  signal blk00000003_sig00000918 : STD_LOGIC; 
  signal blk00000003_sig00000917 : STD_LOGIC; 
  signal blk00000003_sig00000916 : STD_LOGIC; 
  signal blk00000003_sig00000915 : STD_LOGIC; 
  signal blk00000003_sig00000914 : STD_LOGIC; 
  signal blk00000003_sig00000913 : STD_LOGIC; 
  signal blk00000003_sig00000912 : STD_LOGIC; 
  signal blk00000003_sig00000911 : STD_LOGIC; 
  signal blk00000003_sig00000910 : STD_LOGIC; 
  signal blk00000003_sig0000090f : STD_LOGIC; 
  signal blk00000003_sig0000090e : STD_LOGIC; 
  signal blk00000003_sig0000090d : STD_LOGIC; 
  signal blk00000003_sig0000090c : STD_LOGIC; 
  signal blk00000003_sig0000090b : STD_LOGIC; 
  signal blk00000003_sig0000090a : STD_LOGIC; 
  signal blk00000003_sig00000909 : STD_LOGIC; 
  signal blk00000003_sig00000908 : STD_LOGIC; 
  signal blk00000003_sig00000907 : STD_LOGIC; 
  signal blk00000003_sig00000906 : STD_LOGIC; 
  signal blk00000003_sig00000905 : STD_LOGIC; 
  signal blk00000003_sig00000904 : STD_LOGIC; 
  signal blk00000003_sig00000903 : STD_LOGIC; 
  signal blk00000003_sig00000902 : STD_LOGIC; 
  signal blk00000003_sig00000901 : STD_LOGIC; 
  signal blk00000003_sig00000900 : STD_LOGIC; 
  signal blk00000003_sig000008ff : STD_LOGIC; 
  signal blk00000003_sig000008fe : STD_LOGIC; 
  signal blk00000003_sig000008fd : STD_LOGIC; 
  signal blk00000003_sig000008fc : STD_LOGIC; 
  signal blk00000003_sig000008fb : STD_LOGIC; 
  signal blk00000003_sig000008fa : STD_LOGIC; 
  signal blk00000003_sig000008f9 : STD_LOGIC; 
  signal blk00000003_sig000008f8 : STD_LOGIC; 
  signal blk00000003_sig000008f7 : STD_LOGIC; 
  signal blk00000003_sig000008f6 : STD_LOGIC; 
  signal blk00000003_sig000008f5 : STD_LOGIC; 
  signal blk00000003_sig000008f4 : STD_LOGIC; 
  signal blk00000003_sig000008f3 : STD_LOGIC; 
  signal blk00000003_sig000008f2 : STD_LOGIC; 
  signal blk00000003_sig000008f1 : STD_LOGIC; 
  signal blk00000003_sig000008f0 : STD_LOGIC; 
  signal blk00000003_sig000008ef : STD_LOGIC; 
  signal blk00000003_sig000008ee : STD_LOGIC; 
  signal blk00000003_sig000008ed : STD_LOGIC; 
  signal blk00000003_sig000008ec : STD_LOGIC; 
  signal blk00000003_sig000008eb : STD_LOGIC; 
  signal blk00000003_sig000008ea : STD_LOGIC; 
  signal blk00000003_sig000008e9 : STD_LOGIC; 
  signal blk00000003_sig000008e8 : STD_LOGIC; 
  signal blk00000003_sig000008e7 : STD_LOGIC; 
  signal blk00000003_sig000008e6 : STD_LOGIC; 
  signal blk00000003_sig000008e5 : STD_LOGIC; 
  signal blk00000003_sig000008e4 : STD_LOGIC; 
  signal blk00000003_sig000008e3 : STD_LOGIC; 
  signal blk00000003_sig000008e2 : STD_LOGIC; 
  signal blk00000003_sig000008e1 : STD_LOGIC; 
  signal blk00000003_sig000008e0 : STD_LOGIC; 
  signal blk00000003_sig000008df : STD_LOGIC; 
  signal blk00000003_sig000008de : STD_LOGIC; 
  signal blk00000003_sig000008dd : STD_LOGIC; 
  signal blk00000003_sig000008dc : STD_LOGIC; 
  signal blk00000003_sig000008db : STD_LOGIC; 
  signal blk00000003_sig000008da : STD_LOGIC; 
  signal blk00000003_sig000008d9 : STD_LOGIC; 
  signal blk00000003_sig000008d8 : STD_LOGIC; 
  signal blk00000003_sig000008d7 : STD_LOGIC; 
  signal blk00000003_sig000008d6 : STD_LOGIC; 
  signal blk00000003_sig000008d5 : STD_LOGIC; 
  signal blk00000003_sig000008d4 : STD_LOGIC; 
  signal blk00000003_sig000008d3 : STD_LOGIC; 
  signal blk00000003_sig000008d2 : STD_LOGIC; 
  signal blk00000003_sig000008d1 : STD_LOGIC; 
  signal blk00000003_sig000008d0 : STD_LOGIC; 
  signal blk00000003_sig000008cf : STD_LOGIC; 
  signal blk00000003_sig000008ce : STD_LOGIC; 
  signal blk00000003_sig000008cd : STD_LOGIC; 
  signal blk00000003_sig000008cc : STD_LOGIC; 
  signal blk00000003_sig000008cb : STD_LOGIC; 
  signal blk00000003_sig000008ca : STD_LOGIC; 
  signal blk00000003_sig000008c9 : STD_LOGIC; 
  signal blk00000003_sig000008c8 : STD_LOGIC; 
  signal blk00000003_sig000008c7 : STD_LOGIC; 
  signal blk00000003_sig000008c6 : STD_LOGIC; 
  signal blk00000003_sig000008c5 : STD_LOGIC; 
  signal blk00000003_sig000008c4 : STD_LOGIC; 
  signal blk00000003_sig000008c3 : STD_LOGIC; 
  signal blk00000003_sig000008c2 : STD_LOGIC; 
  signal blk00000003_sig000008c1 : STD_LOGIC; 
  signal blk00000003_sig000008c0 : STD_LOGIC; 
  signal blk00000003_sig000008bf : STD_LOGIC; 
  signal blk00000003_sig000008be : STD_LOGIC; 
  signal blk00000003_sig000008bd : STD_LOGIC; 
  signal blk00000003_sig000008bc : STD_LOGIC; 
  signal blk00000003_sig000008bb : STD_LOGIC; 
  signal blk00000003_sig000008ba : STD_LOGIC; 
  signal blk00000003_sig000008b9 : STD_LOGIC; 
  signal blk00000003_sig000008b8 : STD_LOGIC; 
  signal blk00000003_sig000008b7 : STD_LOGIC; 
  signal blk00000003_sig000008b6 : STD_LOGIC; 
  signal blk00000003_sig000008b5 : STD_LOGIC; 
  signal blk00000003_sig000008b4 : STD_LOGIC; 
  signal blk00000003_sig000008b3 : STD_LOGIC; 
  signal blk00000003_sig000008b2 : STD_LOGIC; 
  signal blk00000003_sig000008b1 : STD_LOGIC; 
  signal blk00000003_sig000008b0 : STD_LOGIC; 
  signal blk00000003_sig000008af : STD_LOGIC; 
  signal blk00000003_sig000008ae : STD_LOGIC; 
  signal blk00000003_sig000008ad : STD_LOGIC; 
  signal blk00000003_sig000008ac : STD_LOGIC; 
  signal blk00000003_sig000008ab : STD_LOGIC; 
  signal blk00000003_sig000008aa : STD_LOGIC; 
  signal blk00000003_sig000008a9 : STD_LOGIC; 
  signal blk00000003_sig000008a8 : STD_LOGIC; 
  signal blk00000003_sig000008a7 : STD_LOGIC; 
  signal blk00000003_sig000008a6 : STD_LOGIC; 
  signal blk00000003_sig000008a5 : STD_LOGIC; 
  signal blk00000003_sig000008a4 : STD_LOGIC; 
  signal blk00000003_sig000008a3 : STD_LOGIC; 
  signal blk00000003_sig000008a2 : STD_LOGIC; 
  signal blk00000003_sig000008a1 : STD_LOGIC; 
  signal blk00000003_sig000008a0 : STD_LOGIC; 
  signal blk00000003_sig0000089f : STD_LOGIC; 
  signal blk00000003_sig0000089e : STD_LOGIC; 
  signal blk00000003_sig0000089d : STD_LOGIC; 
  signal blk00000003_sig0000089c : STD_LOGIC; 
  signal blk00000003_sig0000089b : STD_LOGIC; 
  signal blk00000003_sig0000089a : STD_LOGIC; 
  signal blk00000003_sig00000899 : STD_LOGIC; 
  signal blk00000003_sig00000898 : STD_LOGIC; 
  signal blk00000003_sig00000897 : STD_LOGIC; 
  signal blk00000003_sig00000896 : STD_LOGIC; 
  signal blk00000003_sig00000895 : STD_LOGIC; 
  signal blk00000003_sig00000894 : STD_LOGIC; 
  signal blk00000003_sig00000893 : STD_LOGIC; 
  signal blk00000003_sig00000892 : STD_LOGIC; 
  signal blk00000003_sig00000891 : STD_LOGIC; 
  signal blk00000003_sig00000890 : STD_LOGIC; 
  signal blk00000003_sig0000088f : STD_LOGIC; 
  signal blk00000003_sig0000088e : STD_LOGIC; 
  signal blk00000003_sig0000088d : STD_LOGIC; 
  signal blk00000003_sig0000088c : STD_LOGIC; 
  signal blk00000003_sig0000088b : STD_LOGIC; 
  signal blk00000003_sig0000088a : STD_LOGIC; 
  signal blk00000003_sig00000889 : STD_LOGIC; 
  signal blk00000003_sig00000888 : STD_LOGIC; 
  signal blk00000003_sig00000887 : STD_LOGIC; 
  signal blk00000003_sig00000886 : STD_LOGIC; 
  signal blk00000003_sig00000885 : STD_LOGIC; 
  signal blk00000003_sig00000884 : STD_LOGIC; 
  signal blk00000003_sig00000883 : STD_LOGIC; 
  signal blk00000003_sig00000882 : STD_LOGIC; 
  signal blk00000003_sig00000881 : STD_LOGIC; 
  signal blk00000003_sig00000880 : STD_LOGIC; 
  signal blk00000003_sig0000087f : STD_LOGIC; 
  signal blk00000003_sig0000087e : STD_LOGIC; 
  signal blk00000003_sig0000087d : STD_LOGIC; 
  signal blk00000003_sig0000087c : STD_LOGIC; 
  signal blk00000003_sig0000087b : STD_LOGIC; 
  signal blk00000003_sig0000087a : STD_LOGIC; 
  signal blk00000003_sig00000879 : STD_LOGIC; 
  signal blk00000003_sig00000878 : STD_LOGIC; 
  signal blk00000003_sig00000877 : STD_LOGIC; 
  signal blk00000003_sig00000876 : STD_LOGIC; 
  signal blk00000003_sig00000875 : STD_LOGIC; 
  signal blk00000003_sig00000874 : STD_LOGIC; 
  signal blk00000003_sig00000873 : STD_LOGIC; 
  signal blk00000003_sig00000872 : STD_LOGIC; 
  signal blk00000003_sig00000871 : STD_LOGIC; 
  signal blk00000003_sig00000870 : STD_LOGIC; 
  signal blk00000003_sig0000086f : STD_LOGIC; 
  signal blk00000003_sig0000086e : STD_LOGIC; 
  signal blk00000003_sig0000086d : STD_LOGIC; 
  signal blk00000003_sig0000086c : STD_LOGIC; 
  signal blk00000003_sig0000086b : STD_LOGIC; 
  signal blk00000003_sig0000086a : STD_LOGIC; 
  signal blk00000003_sig00000869 : STD_LOGIC; 
  signal blk00000003_sig00000868 : STD_LOGIC; 
  signal blk00000003_sig00000867 : STD_LOGIC; 
  signal blk00000003_sig00000866 : STD_LOGIC; 
  signal blk00000003_sig00000865 : STD_LOGIC; 
  signal blk00000003_sig00000864 : STD_LOGIC; 
  signal blk00000003_sig00000863 : STD_LOGIC; 
  signal blk00000003_sig00000862 : STD_LOGIC; 
  signal blk00000003_sig00000861 : STD_LOGIC; 
  signal blk00000003_sig00000860 : STD_LOGIC; 
  signal blk00000003_sig0000085f : STD_LOGIC; 
  signal blk00000003_sig0000085e : STD_LOGIC; 
  signal blk00000003_sig0000085d : STD_LOGIC; 
  signal blk00000003_sig0000085c : STD_LOGIC; 
  signal blk00000003_sig0000085b : STD_LOGIC; 
  signal blk00000003_sig0000085a : STD_LOGIC; 
  signal blk00000003_sig00000859 : STD_LOGIC; 
  signal blk00000003_sig00000858 : STD_LOGIC; 
  signal blk00000003_sig00000857 : STD_LOGIC; 
  signal blk00000003_sig00000856 : STD_LOGIC; 
  signal blk00000003_sig00000855 : STD_LOGIC; 
  signal blk00000003_sig00000854 : STD_LOGIC; 
  signal blk00000003_sig00000853 : STD_LOGIC; 
  signal blk00000003_sig00000852 : STD_LOGIC; 
  signal blk00000003_sig00000851 : STD_LOGIC; 
  signal blk00000003_sig00000850 : STD_LOGIC; 
  signal blk00000003_sig0000084f : STD_LOGIC; 
  signal blk00000003_sig0000084e : STD_LOGIC; 
  signal blk00000003_sig0000084d : STD_LOGIC; 
  signal blk00000003_sig0000084c : STD_LOGIC; 
  signal blk00000003_sig0000084b : STD_LOGIC; 
  signal blk00000003_sig0000084a : STD_LOGIC; 
  signal blk00000003_sig00000849 : STD_LOGIC; 
  signal blk00000003_sig00000848 : STD_LOGIC; 
  signal blk00000003_sig00000847 : STD_LOGIC; 
  signal blk00000003_sig00000846 : STD_LOGIC; 
  signal blk00000003_sig00000845 : STD_LOGIC; 
  signal blk00000003_sig00000844 : STD_LOGIC; 
  signal blk00000003_sig00000843 : STD_LOGIC; 
  signal blk00000003_sig00000842 : STD_LOGIC; 
  signal blk00000003_sig00000841 : STD_LOGIC; 
  signal blk00000003_sig00000840 : STD_LOGIC; 
  signal blk00000003_sig0000083f : STD_LOGIC; 
  signal blk00000003_sig0000083e : STD_LOGIC; 
  signal blk00000003_sig0000083d : STD_LOGIC; 
  signal blk00000003_sig0000083c : STD_LOGIC; 
  signal blk00000003_sig0000083b : STD_LOGIC; 
  signal blk00000003_sig0000083a : STD_LOGIC; 
  signal blk00000003_sig00000839 : STD_LOGIC; 
  signal blk00000003_sig00000838 : STD_LOGIC; 
  signal blk00000003_sig00000837 : STD_LOGIC; 
  signal blk00000003_sig00000836 : STD_LOGIC; 
  signal blk00000003_sig00000835 : STD_LOGIC; 
  signal blk00000003_sig00000834 : STD_LOGIC; 
  signal blk00000003_sig00000833 : STD_LOGIC; 
  signal blk00000003_sig00000832 : STD_LOGIC; 
  signal blk00000003_sig00000831 : STD_LOGIC; 
  signal blk00000003_sig00000830 : STD_LOGIC; 
  signal blk00000003_sig0000082f : STD_LOGIC; 
  signal blk00000003_sig0000082e : STD_LOGIC; 
  signal blk00000003_sig0000082d : STD_LOGIC; 
  signal blk00000003_sig0000082c : STD_LOGIC; 
  signal blk00000003_sig0000082b : STD_LOGIC; 
  signal blk00000003_sig0000082a : STD_LOGIC; 
  signal blk00000003_sig00000829 : STD_LOGIC; 
  signal blk00000003_sig00000828 : STD_LOGIC; 
  signal blk00000003_sig00000827 : STD_LOGIC; 
  signal blk00000003_sig00000826 : STD_LOGIC; 
  signal blk00000003_sig00000825 : STD_LOGIC; 
  signal blk00000003_sig00000824 : STD_LOGIC; 
  signal blk00000003_sig00000823 : STD_LOGIC; 
  signal blk00000003_sig00000822 : STD_LOGIC; 
  signal blk00000003_sig00000821 : STD_LOGIC; 
  signal blk00000003_sig00000820 : STD_LOGIC; 
  signal blk00000003_sig0000081f : STD_LOGIC; 
  signal blk00000003_sig0000081e : STD_LOGIC; 
  signal blk00000003_sig0000081d : STD_LOGIC; 
  signal blk00000003_sig0000081c : STD_LOGIC; 
  signal blk00000003_sig0000081b : STD_LOGIC; 
  signal blk00000003_sig0000081a : STD_LOGIC; 
  signal blk00000003_sig00000819 : STD_LOGIC; 
  signal blk00000003_sig00000818 : STD_LOGIC; 
  signal blk00000003_sig00000817 : STD_LOGIC; 
  signal blk00000003_sig00000816 : STD_LOGIC; 
  signal blk00000003_sig00000815 : STD_LOGIC; 
  signal blk00000003_sig00000814 : STD_LOGIC; 
  signal blk00000003_sig00000813 : STD_LOGIC; 
  signal blk00000003_sig00000812 : STD_LOGIC; 
  signal blk00000003_sig00000811 : STD_LOGIC; 
  signal blk00000003_sig00000810 : STD_LOGIC; 
  signal blk00000003_sig0000080f : STD_LOGIC; 
  signal blk00000003_sig0000080e : STD_LOGIC; 
  signal blk00000003_sig0000080d : STD_LOGIC; 
  signal blk00000003_sig0000080c : STD_LOGIC; 
  signal blk00000003_sig0000080b : STD_LOGIC; 
  signal blk00000003_sig0000080a : STD_LOGIC; 
  signal blk00000003_sig00000809 : STD_LOGIC; 
  signal blk00000003_sig00000808 : STD_LOGIC; 
  signal blk00000003_sig00000807 : STD_LOGIC; 
  signal blk00000003_sig00000806 : STD_LOGIC; 
  signal blk00000003_sig00000805 : STD_LOGIC; 
  signal blk00000003_sig00000804 : STD_LOGIC; 
  signal blk00000003_sig00000803 : STD_LOGIC; 
  signal blk00000003_sig00000802 : STD_LOGIC; 
  signal blk00000003_sig00000801 : STD_LOGIC; 
  signal blk00000003_sig00000800 : STD_LOGIC; 
  signal blk00000003_sig000007ff : STD_LOGIC; 
  signal blk00000003_sig000007fe : STD_LOGIC; 
  signal blk00000003_sig000007fd : STD_LOGIC; 
  signal blk00000003_sig000007fc : STD_LOGIC; 
  signal blk00000003_sig000007fb : STD_LOGIC; 
  signal blk00000003_sig000007fa : STD_LOGIC; 
  signal blk00000003_sig000007f9 : STD_LOGIC; 
  signal blk00000003_sig000007f8 : STD_LOGIC; 
  signal blk00000003_sig000007f7 : STD_LOGIC; 
  signal blk00000003_sig000007f6 : STD_LOGIC; 
  signal blk00000003_sig000007f5 : STD_LOGIC; 
  signal blk00000003_sig000007f4 : STD_LOGIC; 
  signal blk00000003_sig000007f3 : STD_LOGIC; 
  signal blk00000003_sig000007f2 : STD_LOGIC; 
  signal blk00000003_sig000007f1 : STD_LOGIC; 
  signal blk00000003_sig000007f0 : STD_LOGIC; 
  signal blk00000003_sig000007ef : STD_LOGIC; 
  signal blk00000003_sig000007ee : STD_LOGIC; 
  signal blk00000003_sig000007ed : STD_LOGIC; 
  signal blk00000003_sig000007ec : STD_LOGIC; 
  signal blk00000003_sig000007eb : STD_LOGIC; 
  signal blk00000003_sig000007ea : STD_LOGIC; 
  signal blk00000003_sig000007e9 : STD_LOGIC; 
  signal blk00000003_sig000007e8 : STD_LOGIC; 
  signal blk00000003_sig000007e7 : STD_LOGIC; 
  signal blk00000003_sig000007e6 : STD_LOGIC; 
  signal blk00000003_sig000007e5 : STD_LOGIC; 
  signal blk00000003_sig000007e4 : STD_LOGIC; 
  signal blk00000003_sig000007e3 : STD_LOGIC; 
  signal blk00000003_sig000007e2 : STD_LOGIC; 
  signal blk00000003_sig000007e1 : STD_LOGIC; 
  signal blk00000003_sig000007e0 : STD_LOGIC; 
  signal blk00000003_sig000007df : STD_LOGIC; 
  signal blk00000003_sig000007de : STD_LOGIC; 
  signal blk00000003_sig000007dd : STD_LOGIC; 
  signal blk00000003_sig000007dc : STD_LOGIC; 
  signal blk00000003_sig000007db : STD_LOGIC; 
  signal blk00000003_sig000007da : STD_LOGIC; 
  signal blk00000003_sig000007d9 : STD_LOGIC; 
  signal blk00000003_sig000007d8 : STD_LOGIC; 
  signal blk00000003_sig000007d7 : STD_LOGIC; 
  signal blk00000003_sig000007d6 : STD_LOGIC; 
  signal blk00000003_sig000007d5 : STD_LOGIC; 
  signal blk00000003_sig000007d4 : STD_LOGIC; 
  signal blk00000003_sig000007d3 : STD_LOGIC; 
  signal blk00000003_sig000007d2 : STD_LOGIC; 
  signal blk00000003_sig000007d1 : STD_LOGIC; 
  signal blk00000003_sig000007d0 : STD_LOGIC; 
  signal blk00000003_sig000007cf : STD_LOGIC; 
  signal blk00000003_sig000007ce : STD_LOGIC; 
  signal blk00000003_sig000007cd : STD_LOGIC; 
  signal blk00000003_sig000007cc : STD_LOGIC; 
  signal blk00000003_sig000007cb : STD_LOGIC; 
  signal blk00000003_sig000007ca : STD_LOGIC; 
  signal blk00000003_sig000007c9 : STD_LOGIC; 
  signal blk00000003_sig000007c8 : STD_LOGIC; 
  signal blk00000003_sig000007c7 : STD_LOGIC; 
  signal blk00000003_sig000007c6 : STD_LOGIC; 
  signal blk00000003_sig000007c5 : STD_LOGIC; 
  signal blk00000003_sig000007c4 : STD_LOGIC; 
  signal blk00000003_sig000007c3 : STD_LOGIC; 
  signal blk00000003_sig000007c2 : STD_LOGIC; 
  signal blk00000003_sig000007c1 : STD_LOGIC; 
  signal blk00000003_sig000007c0 : STD_LOGIC; 
  signal blk00000003_sig000007bf : STD_LOGIC; 
  signal blk00000003_sig000007be : STD_LOGIC; 
  signal blk00000003_sig000007bd : STD_LOGIC; 
  signal blk00000003_sig000007bc : STD_LOGIC; 
  signal blk00000003_sig000007bb : STD_LOGIC; 
  signal blk00000003_sig000007ba : STD_LOGIC; 
  signal blk00000003_sig000007b9 : STD_LOGIC; 
  signal blk00000003_sig000007b8 : STD_LOGIC; 
  signal blk00000003_sig000007b7 : STD_LOGIC; 
  signal blk00000003_sig000007b6 : STD_LOGIC; 
  signal blk00000003_sig000007b5 : STD_LOGIC; 
  signal blk00000003_sig000007b4 : STD_LOGIC; 
  signal blk00000003_sig000007b3 : STD_LOGIC; 
  signal blk00000003_sig000007b2 : STD_LOGIC; 
  signal blk00000003_sig000007b1 : STD_LOGIC; 
  signal blk00000003_sig000007b0 : STD_LOGIC; 
  signal blk00000003_sig000007af : STD_LOGIC; 
  signal blk00000003_sig000007ae : STD_LOGIC; 
  signal blk00000003_sig000007ad : STD_LOGIC; 
  signal blk00000003_sig000007ac : STD_LOGIC; 
  signal blk00000003_sig000007ab : STD_LOGIC; 
  signal blk00000003_sig000007aa : STD_LOGIC; 
  signal blk00000003_sig000007a9 : STD_LOGIC; 
  signal blk00000003_sig000007a8 : STD_LOGIC; 
  signal blk00000003_sig000007a7 : STD_LOGIC; 
  signal blk00000003_sig000007a6 : STD_LOGIC; 
  signal blk00000003_sig000007a5 : STD_LOGIC; 
  signal blk00000003_sig000007a4 : STD_LOGIC; 
  signal blk00000003_sig000007a3 : STD_LOGIC; 
  signal blk00000003_sig000007a2 : STD_LOGIC; 
  signal blk00000003_sig000007a1 : STD_LOGIC; 
  signal blk00000003_sig000007a0 : STD_LOGIC; 
  signal blk00000003_sig0000079f : STD_LOGIC; 
  signal blk00000003_sig0000079e : STD_LOGIC; 
  signal blk00000003_sig0000079d : STD_LOGIC; 
  signal blk00000003_sig0000079c : STD_LOGIC; 
  signal blk00000003_sig0000079b : STD_LOGIC; 
  signal blk00000003_sig0000079a : STD_LOGIC; 
  signal blk00000003_sig00000799 : STD_LOGIC; 
  signal blk00000003_sig00000798 : STD_LOGIC; 
  signal blk00000003_sig00000797 : STD_LOGIC; 
  signal blk00000003_sig00000796 : STD_LOGIC; 
  signal blk00000003_sig00000795 : STD_LOGIC; 
  signal blk00000003_sig00000794 : STD_LOGIC; 
  signal blk00000003_sig00000793 : STD_LOGIC; 
  signal blk00000003_sig00000792 : STD_LOGIC; 
  signal blk00000003_sig00000791 : STD_LOGIC; 
  signal blk00000003_sig00000790 : STD_LOGIC; 
  signal blk00000003_sig0000078f : STD_LOGIC; 
  signal blk00000003_sig0000078e : STD_LOGIC; 
  signal blk00000003_sig0000078d : STD_LOGIC; 
  signal blk00000003_sig0000078c : STD_LOGIC; 
  signal blk00000003_sig0000078b : STD_LOGIC; 
  signal blk00000003_sig0000078a : STD_LOGIC; 
  signal blk00000003_sig00000789 : STD_LOGIC; 
  signal blk00000003_sig00000788 : STD_LOGIC; 
  signal blk00000003_sig00000787 : STD_LOGIC; 
  signal blk00000003_sig00000786 : STD_LOGIC; 
  signal blk00000003_sig00000785 : STD_LOGIC; 
  signal blk00000003_sig00000784 : STD_LOGIC; 
  signal blk00000003_sig00000783 : STD_LOGIC; 
  signal blk00000003_sig00000782 : STD_LOGIC; 
  signal blk00000003_sig00000781 : STD_LOGIC; 
  signal blk00000003_sig00000780 : STD_LOGIC; 
  signal blk00000003_sig0000077f : STD_LOGIC; 
  signal blk00000003_sig0000077e : STD_LOGIC; 
  signal blk00000003_sig0000077d : STD_LOGIC; 
  signal blk00000003_sig0000077c : STD_LOGIC; 
  signal blk00000003_sig0000077b : STD_LOGIC; 
  signal blk00000003_sig0000077a : STD_LOGIC; 
  signal blk00000003_sig00000779 : STD_LOGIC; 
  signal blk00000003_sig00000778 : STD_LOGIC; 
  signal blk00000003_sig00000777 : STD_LOGIC; 
  signal blk00000003_sig00000776 : STD_LOGIC; 
  signal blk00000003_sig00000775 : STD_LOGIC; 
  signal blk00000003_sig00000774 : STD_LOGIC; 
  signal blk00000003_sig00000773 : STD_LOGIC; 
  signal blk00000003_sig00000772 : STD_LOGIC; 
  signal blk00000003_sig00000771 : STD_LOGIC; 
  signal blk00000003_sig00000770 : STD_LOGIC; 
  signal blk00000003_sig0000076f : STD_LOGIC; 
  signal blk00000003_sig0000076e : STD_LOGIC; 
  signal blk00000003_sig0000076d : STD_LOGIC; 
  signal blk00000003_sig0000076c : STD_LOGIC; 
  signal blk00000003_sig0000076b : STD_LOGIC; 
  signal blk00000003_sig0000076a : STD_LOGIC; 
  signal blk00000003_sig00000769 : STD_LOGIC; 
  signal blk00000003_sig00000768 : STD_LOGIC; 
  signal blk00000003_sig00000767 : STD_LOGIC; 
  signal blk00000003_sig00000766 : STD_LOGIC; 
  signal blk00000003_sig00000765 : STD_LOGIC; 
  signal blk00000003_sig00000764 : STD_LOGIC; 
  signal blk00000003_sig00000763 : STD_LOGIC; 
  signal blk00000003_sig00000762 : STD_LOGIC; 
  signal blk00000003_sig00000761 : STD_LOGIC; 
  signal blk00000003_sig00000760 : STD_LOGIC; 
  signal blk00000003_sig0000075f : STD_LOGIC; 
  signal blk00000003_sig0000075e : STD_LOGIC; 
  signal blk00000003_sig0000075d : STD_LOGIC; 
  signal blk00000003_sig0000075c : STD_LOGIC; 
  signal blk00000003_sig0000075b : STD_LOGIC; 
  signal blk00000003_sig0000075a : STD_LOGIC; 
  signal blk00000003_sig00000759 : STD_LOGIC; 
  signal blk00000003_sig00000758 : STD_LOGIC; 
  signal blk00000003_sig00000757 : STD_LOGIC; 
  signal blk00000003_sig00000756 : STD_LOGIC; 
  signal blk00000003_sig00000755 : STD_LOGIC; 
  signal blk00000003_sig00000754 : STD_LOGIC; 
  signal blk00000003_sig00000753 : STD_LOGIC; 
  signal blk00000003_sig00000752 : STD_LOGIC; 
  signal blk00000003_sig00000751 : STD_LOGIC; 
  signal blk00000003_sig00000750 : STD_LOGIC; 
  signal blk00000003_sig0000074f : STD_LOGIC; 
  signal blk00000003_sig0000074e : STD_LOGIC; 
  signal blk00000003_sig0000074d : STD_LOGIC; 
  signal blk00000003_sig0000074c : STD_LOGIC; 
  signal blk00000003_sig0000074b : STD_LOGIC; 
  signal blk00000003_sig0000074a : STD_LOGIC; 
  signal blk00000003_sig00000749 : STD_LOGIC; 
  signal blk00000003_sig00000748 : STD_LOGIC; 
  signal blk00000003_sig00000747 : STD_LOGIC; 
  signal blk00000003_sig00000746 : STD_LOGIC; 
  signal blk00000003_sig00000745 : STD_LOGIC; 
  signal blk00000003_sig00000744 : STD_LOGIC; 
  signal blk00000003_sig00000743 : STD_LOGIC; 
  signal blk00000003_sig00000742 : STD_LOGIC; 
  signal blk00000003_sig00000741 : STD_LOGIC; 
  signal blk00000003_sig00000740 : STD_LOGIC; 
  signal blk00000003_sig0000073f : STD_LOGIC; 
  signal blk00000003_sig0000073e : STD_LOGIC; 
  signal blk00000003_sig0000073d : STD_LOGIC; 
  signal blk00000003_sig0000073c : STD_LOGIC; 
  signal blk00000003_sig0000073b : STD_LOGIC; 
  signal blk00000003_sig0000073a : STD_LOGIC; 
  signal blk00000003_sig00000739 : STD_LOGIC; 
  signal blk00000003_sig00000738 : STD_LOGIC; 
  signal blk00000003_sig00000737 : STD_LOGIC; 
  signal blk00000003_sig00000736 : STD_LOGIC; 
  signal blk00000003_sig00000735 : STD_LOGIC; 
  signal blk00000003_sig00000734 : STD_LOGIC; 
  signal blk00000003_sig00000733 : STD_LOGIC; 
  signal blk00000003_sig00000732 : STD_LOGIC; 
  signal blk00000003_sig00000731 : STD_LOGIC; 
  signal blk00000003_sig00000730 : STD_LOGIC; 
  signal blk00000003_sig0000072f : STD_LOGIC; 
  signal blk00000003_sig0000072e : STD_LOGIC; 
  signal blk00000003_sig0000072d : STD_LOGIC; 
  signal blk00000003_sig0000072c : STD_LOGIC; 
  signal blk00000003_sig0000072b : STD_LOGIC; 
  signal blk00000003_sig0000072a : STD_LOGIC; 
  signal blk00000003_sig00000729 : STD_LOGIC; 
  signal blk00000003_sig00000728 : STD_LOGIC; 
  signal blk00000003_sig00000727 : STD_LOGIC; 
  signal blk00000003_sig00000726 : STD_LOGIC; 
  signal blk00000003_sig00000725 : STD_LOGIC; 
  signal blk00000003_sig00000724 : STD_LOGIC; 
  signal blk00000003_sig00000723 : STD_LOGIC; 
  signal blk00000003_sig00000722 : STD_LOGIC; 
  signal blk00000003_sig00000721 : STD_LOGIC; 
  signal blk00000003_sig00000720 : STD_LOGIC; 
  signal blk00000003_sig0000071f : STD_LOGIC; 
  signal blk00000003_sig0000071e : STD_LOGIC; 
  signal blk00000003_sig0000071d : STD_LOGIC; 
  signal blk00000003_sig0000071c : STD_LOGIC; 
  signal blk00000003_sig0000071b : STD_LOGIC; 
  signal blk00000003_sig0000071a : STD_LOGIC; 
  signal blk00000003_sig00000719 : STD_LOGIC; 
  signal blk00000003_sig00000718 : STD_LOGIC; 
  signal blk00000003_sig00000717 : STD_LOGIC; 
  signal blk00000003_sig00000716 : STD_LOGIC; 
  signal blk00000003_sig00000715 : STD_LOGIC; 
  signal blk00000003_sig00000714 : STD_LOGIC; 
  signal blk00000003_sig00000713 : STD_LOGIC; 
  signal blk00000003_sig00000712 : STD_LOGIC; 
  signal blk00000003_sig00000711 : STD_LOGIC; 
  signal blk00000003_sig00000710 : STD_LOGIC; 
  signal blk00000003_sig0000070f : STD_LOGIC; 
  signal blk00000003_sig0000070e : STD_LOGIC; 
  signal blk00000003_sig0000070d : STD_LOGIC; 
  signal blk00000003_sig0000070c : STD_LOGIC; 
  signal blk00000003_sig0000070b : STD_LOGIC; 
  signal blk00000003_sig0000070a : STD_LOGIC; 
  signal blk00000003_sig00000709 : STD_LOGIC; 
  signal blk00000003_sig00000708 : STD_LOGIC; 
  signal blk00000003_sig00000707 : STD_LOGIC; 
  signal blk00000003_sig00000706 : STD_LOGIC; 
  signal blk00000003_sig00000705 : STD_LOGIC; 
  signal blk00000003_sig00000704 : STD_LOGIC; 
  signal blk00000003_sig00000703 : STD_LOGIC; 
  signal blk00000003_sig00000702 : STD_LOGIC; 
  signal blk00000003_sig00000701 : STD_LOGIC; 
  signal blk00000003_sig00000700 : STD_LOGIC; 
  signal blk00000003_sig000006ff : STD_LOGIC; 
  signal blk00000003_sig000006fe : STD_LOGIC; 
  signal blk00000003_sig000006fd : STD_LOGIC; 
  signal blk00000003_sig000006fc : STD_LOGIC; 
  signal blk00000003_sig000006fb : STD_LOGIC; 
  signal blk00000003_sig000006fa : STD_LOGIC; 
  signal blk00000003_sig000006f9 : STD_LOGIC; 
  signal blk00000003_sig000006f8 : STD_LOGIC; 
  signal blk00000003_sig000006f7 : STD_LOGIC; 
  signal blk00000003_sig000006f6 : STD_LOGIC; 
  signal blk00000003_sig000006f5 : STD_LOGIC; 
  signal blk00000003_sig000006f4 : STD_LOGIC; 
  signal blk00000003_sig000006f3 : STD_LOGIC; 
  signal blk00000003_sig000006f2 : STD_LOGIC; 
  signal blk00000003_sig000006f1 : STD_LOGIC; 
  signal blk00000003_sig000006f0 : STD_LOGIC; 
  signal blk00000003_sig000006ef : STD_LOGIC; 
  signal blk00000003_sig000006ee : STD_LOGIC; 
  signal blk00000003_sig000006ed : STD_LOGIC; 
  signal blk00000003_sig000006ec : STD_LOGIC; 
  signal blk00000003_sig000006eb : STD_LOGIC; 
  signal blk00000003_sig000006ea : STD_LOGIC; 
  signal blk00000003_sig000006e9 : STD_LOGIC; 
  signal blk00000003_sig000006e8 : STD_LOGIC; 
  signal blk00000003_sig000006e7 : STD_LOGIC; 
  signal blk00000003_sig000006e6 : STD_LOGIC; 
  signal blk00000003_sig000006e5 : STD_LOGIC; 
  signal blk00000003_sig000006e4 : STD_LOGIC; 
  signal blk00000003_sig000006e3 : STD_LOGIC; 
  signal blk00000003_sig000006e2 : STD_LOGIC; 
  signal blk00000003_sig000006e1 : STD_LOGIC; 
  signal blk00000003_sig000006e0 : STD_LOGIC; 
  signal blk00000003_sig000006df : STD_LOGIC; 
  signal blk00000003_sig000006de : STD_LOGIC; 
  signal blk00000003_sig000006dd : STD_LOGIC; 
  signal blk00000003_sig000006dc : STD_LOGIC; 
  signal blk00000003_sig000006db : STD_LOGIC; 
  signal blk00000003_sig000006da : STD_LOGIC; 
  signal blk00000003_sig000006d9 : STD_LOGIC; 
  signal blk00000003_sig000006d8 : STD_LOGIC; 
  signal blk00000003_sig000006d7 : STD_LOGIC; 
  signal blk00000003_sig000006d6 : STD_LOGIC; 
  signal blk00000003_sig000006d5 : STD_LOGIC; 
  signal blk00000003_sig000006d4 : STD_LOGIC; 
  signal blk00000003_sig000006d3 : STD_LOGIC; 
  signal blk00000003_sig000006d2 : STD_LOGIC; 
  signal blk00000003_sig000006d1 : STD_LOGIC; 
  signal blk00000003_sig000006d0 : STD_LOGIC; 
  signal blk00000003_sig000006cf : STD_LOGIC; 
  signal blk00000003_sig000006ce : STD_LOGIC; 
  signal blk00000003_sig000006cd : STD_LOGIC; 
  signal blk00000003_sig000006cc : STD_LOGIC; 
  signal blk00000003_sig000006cb : STD_LOGIC; 
  signal blk00000003_sig000006ca : STD_LOGIC; 
  signal blk00000003_sig000006c9 : STD_LOGIC; 
  signal blk00000003_sig000006c8 : STD_LOGIC; 
  signal blk00000003_sig000006c7 : STD_LOGIC; 
  signal blk00000003_sig000006c6 : STD_LOGIC; 
  signal blk00000003_sig000006c5 : STD_LOGIC; 
  signal blk00000003_sig000006c4 : STD_LOGIC; 
  signal blk00000003_sig000006c3 : STD_LOGIC; 
  signal blk00000003_sig000006c2 : STD_LOGIC; 
  signal blk00000003_sig000006c1 : STD_LOGIC; 
  signal blk00000003_sig000006c0 : STD_LOGIC; 
  signal blk00000003_sig000006bf : STD_LOGIC; 
  signal blk00000003_sig000006be : STD_LOGIC; 
  signal blk00000003_sig000006bd : STD_LOGIC; 
  signal blk00000003_sig000006bc : STD_LOGIC; 
  signal blk00000003_sig000006bb : STD_LOGIC; 
  signal blk00000003_sig000006ba : STD_LOGIC; 
  signal blk00000003_sig000006b9 : STD_LOGIC; 
  signal blk00000003_sig000006b8 : STD_LOGIC; 
  signal blk00000003_sig000006b7 : STD_LOGIC; 
  signal blk00000003_sig000006b6 : STD_LOGIC; 
  signal blk00000003_sig000006b5 : STD_LOGIC; 
  signal blk00000003_sig000006b4 : STD_LOGIC; 
  signal blk00000003_sig000006b3 : STD_LOGIC; 
  signal blk00000003_sig000006b2 : STD_LOGIC; 
  signal blk00000003_sig000006b1 : STD_LOGIC; 
  signal blk00000003_sig000006b0 : STD_LOGIC; 
  signal blk00000003_sig000006af : STD_LOGIC; 
  signal blk00000003_sig000006ae : STD_LOGIC; 
  signal blk00000003_sig000006ad : STD_LOGIC; 
  signal blk00000003_sig000006ac : STD_LOGIC; 
  signal blk00000003_sig000006ab : STD_LOGIC; 
  signal blk00000003_sig000006aa : STD_LOGIC; 
  signal blk00000003_sig000006a9 : STD_LOGIC; 
  signal blk00000003_sig000006a8 : STD_LOGIC; 
  signal blk00000003_sig000006a7 : STD_LOGIC; 
  signal blk00000003_sig000006a6 : STD_LOGIC; 
  signal blk00000003_sig000006a5 : STD_LOGIC; 
  signal blk00000003_sig000006a4 : STD_LOGIC; 
  signal blk00000003_sig000006a3 : STD_LOGIC; 
  signal blk00000003_sig000006a2 : STD_LOGIC; 
  signal blk00000003_sig000006a1 : STD_LOGIC; 
  signal blk00000003_sig000006a0 : STD_LOGIC; 
  signal blk00000003_sig0000069f : STD_LOGIC; 
  signal blk00000003_sig0000069e : STD_LOGIC; 
  signal blk00000003_sig0000069d : STD_LOGIC; 
  signal blk00000003_sig0000069c : STD_LOGIC; 
  signal blk00000003_sig0000069b : STD_LOGIC; 
  signal blk00000003_sig0000069a : STD_LOGIC; 
  signal blk00000003_sig00000699 : STD_LOGIC; 
  signal blk00000003_sig00000698 : STD_LOGIC; 
  signal blk00000003_sig00000697 : STD_LOGIC; 
  signal blk00000003_sig00000696 : STD_LOGIC; 
  signal blk00000003_sig00000695 : STD_LOGIC; 
  signal blk00000003_sig00000694 : STD_LOGIC; 
  signal blk00000003_sig00000693 : STD_LOGIC; 
  signal blk00000003_sig00000692 : STD_LOGIC; 
  signal blk00000003_sig00000691 : STD_LOGIC; 
  signal blk00000003_sig00000690 : STD_LOGIC; 
  signal blk00000003_sig0000068f : STD_LOGIC; 
  signal blk00000003_sig0000068e : STD_LOGIC; 
  signal blk00000003_sig0000068d : STD_LOGIC; 
  signal blk00000003_sig0000068c : STD_LOGIC; 
  signal blk00000003_sig0000068b : STD_LOGIC; 
  signal blk00000003_sig0000068a : STD_LOGIC; 
  signal blk00000003_sig00000689 : STD_LOGIC; 
  signal blk00000003_sig00000688 : STD_LOGIC; 
  signal blk00000003_sig00000687 : STD_LOGIC; 
  signal blk00000003_sig00000686 : STD_LOGIC; 
  signal blk00000003_sig00000685 : STD_LOGIC; 
  signal blk00000003_sig00000684 : STD_LOGIC; 
  signal blk00000003_sig00000683 : STD_LOGIC; 
  signal blk00000003_sig00000682 : STD_LOGIC; 
  signal blk00000003_sig00000681 : STD_LOGIC; 
  signal blk00000003_sig00000680 : STD_LOGIC; 
  signal blk00000003_sig0000067f : STD_LOGIC; 
  signal blk00000003_sig0000067e : STD_LOGIC; 
  signal blk00000003_sig0000067d : STD_LOGIC; 
  signal blk00000003_sig0000067c : STD_LOGIC; 
  signal blk00000003_sig0000067b : STD_LOGIC; 
  signal blk00000003_sig0000067a : STD_LOGIC; 
  signal blk00000003_sig00000679 : STD_LOGIC; 
  signal blk00000003_sig00000678 : STD_LOGIC; 
  signal blk00000003_sig00000677 : STD_LOGIC; 
  signal blk00000003_sig00000676 : STD_LOGIC; 
  signal blk00000003_sig00000675 : STD_LOGIC; 
  signal blk00000003_sig00000674 : STD_LOGIC; 
  signal blk00000003_sig00000673 : STD_LOGIC; 
  signal blk00000003_sig00000672 : STD_LOGIC; 
  signal blk00000003_sig00000671 : STD_LOGIC; 
  signal blk00000003_sig00000670 : STD_LOGIC; 
  signal blk00000003_sig0000066f : STD_LOGIC; 
  signal blk00000003_sig0000066e : STD_LOGIC; 
  signal blk00000003_sig0000066d : STD_LOGIC; 
  signal blk00000003_sig0000066c : STD_LOGIC; 
  signal blk00000003_sig0000066b : STD_LOGIC; 
  signal blk00000003_sig0000066a : STD_LOGIC; 
  signal blk00000003_sig00000669 : STD_LOGIC; 
  signal blk00000003_sig00000668 : STD_LOGIC; 
  signal blk00000003_sig00000667 : STD_LOGIC; 
  signal blk00000003_sig00000666 : STD_LOGIC; 
  signal blk00000003_sig00000665 : STD_LOGIC; 
  signal blk00000003_sig00000664 : STD_LOGIC; 
  signal blk00000003_sig00000663 : STD_LOGIC; 
  signal blk00000003_sig00000662 : STD_LOGIC; 
  signal blk00000003_sig00000661 : STD_LOGIC; 
  signal blk00000003_sig00000660 : STD_LOGIC; 
  signal blk00000003_sig0000065f : STD_LOGIC; 
  signal blk00000003_sig0000065e : STD_LOGIC; 
  signal blk00000003_sig0000065d : STD_LOGIC; 
  signal blk00000003_sig0000065c : STD_LOGIC; 
  signal blk00000003_sig0000065b : STD_LOGIC; 
  signal blk00000003_sig0000065a : STD_LOGIC; 
  signal blk00000003_sig00000659 : STD_LOGIC; 
  signal blk00000003_sig00000658 : STD_LOGIC; 
  signal blk00000003_sig00000657 : STD_LOGIC; 
  signal blk00000003_sig00000656 : STD_LOGIC; 
  signal blk00000003_sig00000655 : STD_LOGIC; 
  signal blk00000003_sig00000654 : STD_LOGIC; 
  signal blk00000003_sig00000653 : STD_LOGIC; 
  signal blk00000003_sig00000652 : STD_LOGIC; 
  signal blk00000003_sig00000651 : STD_LOGIC; 
  signal blk00000003_sig00000650 : STD_LOGIC; 
  signal blk00000003_sig0000064f : STD_LOGIC; 
  signal blk00000003_sig0000064e : STD_LOGIC; 
  signal blk00000003_sig0000064d : STD_LOGIC; 
  signal blk00000003_sig0000064c : STD_LOGIC; 
  signal blk00000003_sig0000064b : STD_LOGIC; 
  signal blk00000003_sig0000064a : STD_LOGIC; 
  signal blk00000003_sig00000649 : STD_LOGIC; 
  signal blk00000003_sig00000648 : STD_LOGIC; 
  signal blk00000003_sig00000647 : STD_LOGIC; 
  signal blk00000003_sig00000646 : STD_LOGIC; 
  signal blk00000003_sig00000645 : STD_LOGIC; 
  signal blk00000003_sig00000644 : STD_LOGIC; 
  signal blk00000003_sig00000643 : STD_LOGIC; 
  signal blk00000003_sig00000642 : STD_LOGIC; 
  signal blk00000003_sig00000641 : STD_LOGIC; 
  signal blk00000003_sig00000640 : STD_LOGIC; 
  signal blk00000003_sig0000063f : STD_LOGIC; 
  signal blk00000003_sig0000063e : STD_LOGIC; 
  signal blk00000003_sig0000063d : STD_LOGIC; 
  signal blk00000003_sig0000063c : STD_LOGIC; 
  signal blk00000003_sig0000063b : STD_LOGIC; 
  signal blk00000003_sig0000063a : STD_LOGIC; 
  signal blk00000003_sig00000639 : STD_LOGIC; 
  signal blk00000003_sig00000638 : STD_LOGIC; 
  signal blk00000003_sig00000637 : STD_LOGIC; 
  signal blk00000003_sig00000636 : STD_LOGIC; 
  signal blk00000003_sig00000635 : STD_LOGIC; 
  signal blk00000003_sig00000634 : STD_LOGIC; 
  signal blk00000003_sig00000633 : STD_LOGIC; 
  signal blk00000003_sig00000632 : STD_LOGIC; 
  signal blk00000003_sig00000631 : STD_LOGIC; 
  signal blk00000003_sig00000630 : STD_LOGIC; 
  signal blk00000003_sig0000062f : STD_LOGIC; 
  signal blk00000003_sig0000062e : STD_LOGIC; 
  signal blk00000003_sig0000062d : STD_LOGIC; 
  signal blk00000003_sig0000062c : STD_LOGIC; 
  signal blk00000003_sig0000062b : STD_LOGIC; 
  signal blk00000003_sig0000062a : STD_LOGIC; 
  signal blk00000003_sig00000629 : STD_LOGIC; 
  signal blk00000003_sig00000628 : STD_LOGIC; 
  signal blk00000003_sig00000627 : STD_LOGIC; 
  signal blk00000003_sig00000626 : STD_LOGIC; 
  signal blk00000003_sig00000625 : STD_LOGIC; 
  signal blk00000003_sig00000624 : STD_LOGIC; 
  signal blk00000003_sig00000623 : STD_LOGIC; 
  signal blk00000003_sig00000622 : STD_LOGIC; 
  signal blk00000003_sig00000621 : STD_LOGIC; 
  signal blk00000003_sig00000620 : STD_LOGIC; 
  signal blk00000003_sig0000061f : STD_LOGIC; 
  signal blk00000003_sig0000061e : STD_LOGIC; 
  signal blk00000003_sig0000061d : STD_LOGIC; 
  signal blk00000003_sig0000061c : STD_LOGIC; 
  signal blk00000003_sig0000061b : STD_LOGIC; 
  signal blk00000003_sig0000061a : STD_LOGIC; 
  signal blk00000003_sig00000619 : STD_LOGIC; 
  signal blk00000003_sig00000618 : STD_LOGIC; 
  signal blk00000003_sig00000617 : STD_LOGIC; 
  signal blk00000003_sig00000616 : STD_LOGIC; 
  signal blk00000003_sig00000615 : STD_LOGIC; 
  signal blk00000003_sig00000614 : STD_LOGIC; 
  signal blk00000003_sig00000613 : STD_LOGIC; 
  signal blk00000003_sig00000612 : STD_LOGIC; 
  signal blk00000003_sig00000611 : STD_LOGIC; 
  signal blk00000003_sig00000610 : STD_LOGIC; 
  signal blk00000003_sig0000060f : STD_LOGIC; 
  signal blk00000003_sig0000060e : STD_LOGIC; 
  signal blk00000003_sig0000060d : STD_LOGIC; 
  signal blk00000003_sig0000060c : STD_LOGIC; 
  signal blk00000003_sig0000060b : STD_LOGIC; 
  signal blk00000003_sig0000060a : STD_LOGIC; 
  signal blk00000003_sig00000609 : STD_LOGIC; 
  signal blk00000003_sig00000608 : STD_LOGIC; 
  signal blk00000003_sig00000607 : STD_LOGIC; 
  signal blk00000003_sig00000606 : STD_LOGIC; 
  signal blk00000003_sig00000605 : STD_LOGIC; 
  signal blk00000003_sig00000604 : STD_LOGIC; 
  signal blk00000003_sig00000603 : STD_LOGIC; 
  signal blk00000003_sig00000602 : STD_LOGIC; 
  signal blk00000003_sig00000601 : STD_LOGIC; 
  signal blk00000003_sig00000600 : STD_LOGIC; 
  signal blk00000003_sig000005ff : STD_LOGIC; 
  signal blk00000003_sig000005fe : STD_LOGIC; 
  signal blk00000003_sig000005fd : STD_LOGIC; 
  signal blk00000003_sig000005fc : STD_LOGIC; 
  signal blk00000003_sig000005fb : STD_LOGIC; 
  signal blk00000003_sig000005fa : STD_LOGIC; 
  signal blk00000003_sig000005f9 : STD_LOGIC; 
  signal blk00000003_sig000005f8 : STD_LOGIC; 
  signal blk00000003_sig000005f7 : STD_LOGIC; 
  signal blk00000003_sig000005f6 : STD_LOGIC; 
  signal blk00000003_sig000005f5 : STD_LOGIC; 
  signal blk00000003_sig000005f4 : STD_LOGIC; 
  signal blk00000003_sig000005f3 : STD_LOGIC; 
  signal blk00000003_sig000005f2 : STD_LOGIC; 
  signal blk00000003_sig000005f1 : STD_LOGIC; 
  signal blk00000003_sig000005f0 : STD_LOGIC; 
  signal blk00000003_sig000005ef : STD_LOGIC; 
  signal blk00000003_sig000005ee : STD_LOGIC; 
  signal blk00000003_sig000005ed : STD_LOGIC; 
  signal blk00000003_sig000005ec : STD_LOGIC; 
  signal blk00000003_sig000005eb : STD_LOGIC; 
  signal blk00000003_sig000005ea : STD_LOGIC; 
  signal blk00000003_sig000005e9 : STD_LOGIC; 
  signal blk00000003_sig000005e8 : STD_LOGIC; 
  signal blk00000003_sig000005e7 : STD_LOGIC; 
  signal blk00000003_sig000005e6 : STD_LOGIC; 
  signal blk00000003_sig000005e5 : STD_LOGIC; 
  signal blk00000003_sig000005e4 : STD_LOGIC; 
  signal blk00000003_sig000005e3 : STD_LOGIC; 
  signal blk00000003_sig000005e2 : STD_LOGIC; 
  signal blk00000003_sig000005e1 : STD_LOGIC; 
  signal blk00000003_sig000005e0 : STD_LOGIC; 
  signal blk00000003_sig000005df : STD_LOGIC; 
  signal blk00000003_sig000005de : STD_LOGIC; 
  signal blk00000003_sig000005dd : STD_LOGIC; 
  signal blk00000003_sig000005dc : STD_LOGIC; 
  signal blk00000003_sig000005db : STD_LOGIC; 
  signal blk00000003_sig000005da : STD_LOGIC; 
  signal blk00000003_sig000005d9 : STD_LOGIC; 
  signal blk00000003_sig000005d8 : STD_LOGIC; 
  signal blk00000003_sig000005d7 : STD_LOGIC; 
  signal blk00000003_sig000005d6 : STD_LOGIC; 
  signal blk00000003_sig000005d5 : STD_LOGIC; 
  signal blk00000003_sig000005d4 : STD_LOGIC; 
  signal blk00000003_sig000005d3 : STD_LOGIC; 
  signal blk00000003_sig000005d2 : STD_LOGIC; 
  signal blk00000003_sig000005d1 : STD_LOGIC; 
  signal blk00000003_sig000005d0 : STD_LOGIC; 
  signal blk00000003_sig000005cf : STD_LOGIC; 
  signal blk00000003_sig000005ce : STD_LOGIC; 
  signal blk00000003_sig000005cd : STD_LOGIC; 
  signal blk00000003_sig000005cc : STD_LOGIC; 
  signal blk00000003_sig000005cb : STD_LOGIC; 
  signal blk00000003_sig000005ca : STD_LOGIC; 
  signal blk00000003_sig000005c9 : STD_LOGIC; 
  signal blk00000003_sig000005c8 : STD_LOGIC; 
  signal blk00000003_sig000005c7 : STD_LOGIC; 
  signal blk00000003_sig000005c6 : STD_LOGIC; 
  signal blk00000003_sig000005c5 : STD_LOGIC; 
  signal blk00000003_sig000005c4 : STD_LOGIC; 
  signal blk00000003_sig000005c3 : STD_LOGIC; 
  signal blk00000003_sig000005c2 : STD_LOGIC; 
  signal blk00000003_sig000005c1 : STD_LOGIC; 
  signal blk00000003_sig000005c0 : STD_LOGIC; 
  signal blk00000003_sig000005bf : STD_LOGIC; 
  signal blk00000003_sig000005be : STD_LOGIC; 
  signal blk00000003_sig000005bd : STD_LOGIC; 
  signal blk00000003_sig000005bc : STD_LOGIC; 
  signal blk00000003_sig000005bb : STD_LOGIC; 
  signal blk00000003_sig000005ba : STD_LOGIC; 
  signal blk00000003_sig000005b9 : STD_LOGIC; 
  signal blk00000003_sig000005b8 : STD_LOGIC; 
  signal blk00000003_sig000005b7 : STD_LOGIC; 
  signal blk00000003_sig000005b6 : STD_LOGIC; 
  signal blk00000003_sig000005b5 : STD_LOGIC; 
  signal blk00000003_sig000005b4 : STD_LOGIC; 
  signal blk00000003_sig000005b3 : STD_LOGIC; 
  signal blk00000003_sig000005b2 : STD_LOGIC; 
  signal blk00000003_sig000005b1 : STD_LOGIC; 
  signal blk00000003_sig000005b0 : STD_LOGIC; 
  signal blk00000003_sig000005af : STD_LOGIC; 
  signal blk00000003_sig000005ae : STD_LOGIC; 
  signal blk00000003_sig000005ad : STD_LOGIC; 
  signal blk00000003_sig000005ac : STD_LOGIC; 
  signal blk00000003_sig000005ab : STD_LOGIC; 
  signal blk00000003_sig000005aa : STD_LOGIC; 
  signal blk00000003_sig000005a9 : STD_LOGIC; 
  signal blk00000003_sig000005a8 : STD_LOGIC; 
  signal blk00000003_sig000005a7 : STD_LOGIC; 
  signal blk00000003_sig000005a6 : STD_LOGIC; 
  signal blk00000003_sig000005a5 : STD_LOGIC; 
  signal blk00000003_sig000005a4 : STD_LOGIC; 
  signal blk00000003_sig000005a3 : STD_LOGIC; 
  signal blk00000003_sig000005a2 : STD_LOGIC; 
  signal blk00000003_sig000005a1 : STD_LOGIC; 
  signal blk00000003_sig000005a0 : STD_LOGIC; 
  signal blk00000003_sig0000059f : STD_LOGIC; 
  signal blk00000003_sig0000059e : STD_LOGIC; 
  signal blk00000003_sig0000059d : STD_LOGIC; 
  signal blk00000003_sig0000059c : STD_LOGIC; 
  signal blk00000003_sig0000059b : STD_LOGIC; 
  signal blk00000003_sig0000059a : STD_LOGIC; 
  signal blk00000003_sig00000599 : STD_LOGIC; 
  signal blk00000003_sig00000598 : STD_LOGIC; 
  signal blk00000003_sig00000597 : STD_LOGIC; 
  signal blk00000003_sig00000596 : STD_LOGIC; 
  signal blk00000003_sig00000595 : STD_LOGIC; 
  signal blk00000003_sig00000594 : STD_LOGIC; 
  signal blk00000003_sig00000593 : STD_LOGIC; 
  signal blk00000003_sig00000592 : STD_LOGIC; 
  signal blk00000003_sig00000591 : STD_LOGIC; 
  signal blk00000003_sig00000590 : STD_LOGIC; 
  signal blk00000003_sig0000058f : STD_LOGIC; 
  signal blk00000003_sig0000058e : STD_LOGIC; 
  signal blk00000003_sig0000058d : STD_LOGIC; 
  signal blk00000003_sig0000058c : STD_LOGIC; 
  signal blk00000003_sig0000058b : STD_LOGIC; 
  signal blk00000003_sig0000058a : STD_LOGIC; 
  signal blk00000003_sig00000589 : STD_LOGIC; 
  signal blk00000003_sig00000588 : STD_LOGIC; 
  signal blk00000003_sig00000587 : STD_LOGIC; 
  signal blk00000003_sig00000586 : STD_LOGIC; 
  signal blk00000003_sig00000585 : STD_LOGIC; 
  signal blk00000003_sig00000584 : STD_LOGIC; 
  signal blk00000003_sig00000583 : STD_LOGIC; 
  signal blk00000003_sig00000582 : STD_LOGIC; 
  signal blk00000003_sig00000581 : STD_LOGIC; 
  signal blk00000003_sig00000580 : STD_LOGIC; 
  signal blk00000003_sig0000057f : STD_LOGIC; 
  signal blk00000003_sig0000057e : STD_LOGIC; 
  signal blk00000003_sig0000057d : STD_LOGIC; 
  signal blk00000003_sig0000057c : STD_LOGIC; 
  signal blk00000003_sig0000057b : STD_LOGIC; 
  signal blk00000003_sig0000057a : STD_LOGIC; 
  signal blk00000003_sig00000579 : STD_LOGIC; 
  signal blk00000003_sig00000578 : STD_LOGIC; 
  signal blk00000003_sig00000577 : STD_LOGIC; 
  signal blk00000003_sig00000576 : STD_LOGIC; 
  signal blk00000003_sig00000575 : STD_LOGIC; 
  signal blk00000003_sig00000574 : STD_LOGIC; 
  signal blk00000003_sig00000573 : STD_LOGIC; 
  signal blk00000003_sig00000572 : STD_LOGIC; 
  signal blk00000003_sig00000571 : STD_LOGIC; 
  signal blk00000003_sig00000570 : STD_LOGIC; 
  signal blk00000003_sig0000056f : STD_LOGIC; 
  signal blk00000003_sig0000056e : STD_LOGIC; 
  signal blk00000003_sig0000056d : STD_LOGIC; 
  signal blk00000003_sig0000056c : STD_LOGIC; 
  signal blk00000003_sig0000056b : STD_LOGIC; 
  signal blk00000003_sig0000056a : STD_LOGIC; 
  signal blk00000003_sig00000569 : STD_LOGIC; 
  signal blk00000003_sig00000568 : STD_LOGIC; 
  signal blk00000003_sig00000567 : STD_LOGIC; 
  signal blk00000003_sig00000566 : STD_LOGIC; 
  signal blk00000003_sig00000565 : STD_LOGIC; 
  signal blk00000003_sig00000564 : STD_LOGIC; 
  signal blk00000003_sig00000563 : STD_LOGIC; 
  signal blk00000003_sig00000562 : STD_LOGIC; 
  signal blk00000003_sig00000561 : STD_LOGIC; 
  signal blk00000003_sig00000560 : STD_LOGIC; 
  signal blk00000003_sig0000055f : STD_LOGIC; 
  signal blk00000003_sig0000055e : STD_LOGIC; 
  signal blk00000003_sig0000055d : STD_LOGIC; 
  signal blk00000003_sig0000055c : STD_LOGIC; 
  signal blk00000003_sig0000055b : STD_LOGIC; 
  signal blk00000003_sig0000055a : STD_LOGIC; 
  signal blk00000003_sig00000559 : STD_LOGIC; 
  signal blk00000003_sig00000558 : STD_LOGIC; 
  signal blk00000003_sig00000557 : STD_LOGIC; 
  signal blk00000003_sig00000556 : STD_LOGIC; 
  signal blk00000003_sig00000555 : STD_LOGIC; 
  signal blk00000003_sig00000554 : STD_LOGIC; 
  signal blk00000003_sig00000553 : STD_LOGIC; 
  signal blk00000003_sig00000552 : STD_LOGIC; 
  signal blk00000003_sig00000551 : STD_LOGIC; 
  signal blk00000003_sig00000550 : STD_LOGIC; 
  signal blk00000003_sig0000054f : STD_LOGIC; 
  signal blk00000003_sig0000054e : STD_LOGIC; 
  signal blk00000003_sig0000054d : STD_LOGIC; 
  signal blk00000003_sig0000054c : STD_LOGIC; 
  signal blk00000003_sig0000054b : STD_LOGIC; 
  signal blk00000003_sig0000054a : STD_LOGIC; 
  signal blk00000003_sig00000549 : STD_LOGIC; 
  signal blk00000003_sig00000548 : STD_LOGIC; 
  signal blk00000003_sig00000547 : STD_LOGIC; 
  signal blk00000003_sig00000546 : STD_LOGIC; 
  signal blk00000003_sig00000545 : STD_LOGIC; 
  signal blk00000003_sig00000544 : STD_LOGIC; 
  signal blk00000003_sig00000543 : STD_LOGIC; 
  signal blk00000003_sig00000542 : STD_LOGIC; 
  signal blk00000003_sig00000541 : STD_LOGIC; 
  signal blk00000003_sig00000540 : STD_LOGIC; 
  signal blk00000003_sig0000053f : STD_LOGIC; 
  signal blk00000003_sig0000053e : STD_LOGIC; 
  signal blk00000003_sig0000053d : STD_LOGIC; 
  signal blk00000003_sig0000053c : STD_LOGIC; 
  signal blk00000003_sig0000053b : STD_LOGIC; 
  signal blk00000003_sig0000053a : STD_LOGIC; 
  signal blk00000003_sig00000539 : STD_LOGIC; 
  signal blk00000003_sig00000538 : STD_LOGIC; 
  signal blk00000003_sig00000537 : STD_LOGIC; 
  signal blk00000003_sig00000536 : STD_LOGIC; 
  signal blk00000003_sig00000535 : STD_LOGIC; 
  signal blk00000003_sig00000534 : STD_LOGIC; 
  signal blk00000003_sig00000533 : STD_LOGIC; 
  signal blk00000003_sig00000532 : STD_LOGIC; 
  signal blk00000003_sig00000531 : STD_LOGIC; 
  signal blk00000003_sig00000530 : STD_LOGIC; 
  signal blk00000003_sig0000052f : STD_LOGIC; 
  signal blk00000003_sig0000052e : STD_LOGIC; 
  signal blk00000003_sig0000052d : STD_LOGIC; 
  signal blk00000003_sig0000052c : STD_LOGIC; 
  signal blk00000003_sig0000052b : STD_LOGIC; 
  signal blk00000003_sig0000052a : STD_LOGIC; 
  signal blk00000003_sig00000529 : STD_LOGIC; 
  signal blk00000003_sig00000528 : STD_LOGIC; 
  signal blk00000003_sig00000527 : STD_LOGIC; 
  signal blk00000003_sig00000526 : STD_LOGIC; 
  signal blk00000003_sig00000525 : STD_LOGIC; 
  signal blk00000003_sig00000524 : STD_LOGIC; 
  signal blk00000003_sig00000523 : STD_LOGIC; 
  signal blk00000003_sig00000522 : STD_LOGIC; 
  signal blk00000003_sig00000521 : STD_LOGIC; 
  signal blk00000003_sig00000520 : STD_LOGIC; 
  signal blk00000003_sig0000051f : STD_LOGIC; 
  signal blk00000003_sig0000051e : STD_LOGIC; 
  signal blk00000003_sig0000051d : STD_LOGIC; 
  signal blk00000003_sig0000051c : STD_LOGIC; 
  signal blk00000003_sig0000051b : STD_LOGIC; 
  signal blk00000003_sig0000051a : STD_LOGIC; 
  signal blk00000003_sig00000519 : STD_LOGIC; 
  signal blk00000003_sig00000518 : STD_LOGIC; 
  signal blk00000003_sig00000517 : STD_LOGIC; 
  signal blk00000003_sig00000516 : STD_LOGIC; 
  signal blk00000003_sig00000515 : STD_LOGIC; 
  signal blk00000003_sig00000514 : STD_LOGIC; 
  signal blk00000003_sig00000513 : STD_LOGIC; 
  signal blk00000003_sig00000512 : STD_LOGIC; 
  signal blk00000003_sig00000511 : STD_LOGIC; 
  signal blk00000003_sig00000510 : STD_LOGIC; 
  signal blk00000003_sig0000050f : STD_LOGIC; 
  signal blk00000003_sig0000050e : STD_LOGIC; 
  signal blk00000003_sig0000050d : STD_LOGIC; 
  signal blk00000003_sig0000050c : STD_LOGIC; 
  signal blk00000003_sig0000050b : STD_LOGIC; 
  signal blk00000003_sig0000050a : STD_LOGIC; 
  signal blk00000003_sig00000509 : STD_LOGIC; 
  signal blk00000003_sig00000508 : STD_LOGIC; 
  signal blk00000003_sig00000507 : STD_LOGIC; 
  signal blk00000003_sig00000506 : STD_LOGIC; 
  signal blk00000003_sig00000505 : STD_LOGIC; 
  signal blk00000003_sig00000504 : STD_LOGIC; 
  signal blk00000003_sig00000503 : STD_LOGIC; 
  signal blk00000003_sig00000502 : STD_LOGIC; 
  signal blk00000003_sig00000501 : STD_LOGIC; 
  signal blk00000003_sig00000500 : STD_LOGIC; 
  signal blk00000003_sig000004ff : STD_LOGIC; 
  signal blk00000003_sig000004fe : STD_LOGIC; 
  signal blk00000003_sig000004fd : STD_LOGIC; 
  signal blk00000003_sig000004fc : STD_LOGIC; 
  signal blk00000003_sig000004fb : STD_LOGIC; 
  signal blk00000003_sig000004fa : STD_LOGIC; 
  signal blk00000003_sig000004f9 : STD_LOGIC; 
  signal blk00000003_sig000004f8 : STD_LOGIC; 
  signal blk00000003_sig000004f7 : STD_LOGIC; 
  signal blk00000003_sig000004f6 : STD_LOGIC; 
  signal blk00000003_sig000004f5 : STD_LOGIC; 
  signal blk00000003_sig000004f4 : STD_LOGIC; 
  signal blk00000003_sig000004f3 : STD_LOGIC; 
  signal blk00000003_sig000004f2 : STD_LOGIC; 
  signal blk00000003_sig000004f1 : STD_LOGIC; 
  signal blk00000003_sig000004f0 : STD_LOGIC; 
  signal blk00000003_sig000004ef : STD_LOGIC; 
  signal blk00000003_sig000004ee : STD_LOGIC; 
  signal blk00000003_sig000004ed : STD_LOGIC; 
  signal blk00000003_sig000004ec : STD_LOGIC; 
  signal blk00000003_sig000004eb : STD_LOGIC; 
  signal blk00000003_sig000004ea : STD_LOGIC; 
  signal blk00000003_sig000004e9 : STD_LOGIC; 
  signal blk00000003_sig000004e8 : STD_LOGIC; 
  signal blk00000003_sig000004e7 : STD_LOGIC; 
  signal blk00000003_sig000004e6 : STD_LOGIC; 
  signal blk00000003_sig000004e5 : STD_LOGIC; 
  signal blk00000003_sig000004e4 : STD_LOGIC; 
  signal blk00000003_sig000004e3 : STD_LOGIC; 
  signal blk00000003_sig000004e2 : STD_LOGIC; 
  signal blk00000003_sig000004e1 : STD_LOGIC; 
  signal blk00000003_sig000004e0 : STD_LOGIC; 
  signal blk00000003_sig000004df : STD_LOGIC; 
  signal blk00000003_sig000004de : STD_LOGIC; 
  signal blk00000003_sig000004dd : STD_LOGIC; 
  signal blk00000003_sig000004dc : STD_LOGIC; 
  signal blk00000003_sig000004db : STD_LOGIC; 
  signal blk00000003_sig000004da : STD_LOGIC; 
  signal blk00000003_sig000004d9 : STD_LOGIC; 
  signal blk00000003_sig000004d8 : STD_LOGIC; 
  signal blk00000003_sig000004d7 : STD_LOGIC; 
  signal blk00000003_sig000004d6 : STD_LOGIC; 
  signal blk00000003_sig000004d5 : STD_LOGIC; 
  signal blk00000003_sig000004d4 : STD_LOGIC; 
  signal blk00000003_sig000004d3 : STD_LOGIC; 
  signal blk00000003_sig000004d2 : STD_LOGIC; 
  signal blk00000003_sig000004d1 : STD_LOGIC; 
  signal blk00000003_sig000004d0 : STD_LOGIC; 
  signal blk00000003_sig000004cf : STD_LOGIC; 
  signal blk00000003_sig000004ce : STD_LOGIC; 
  signal blk00000003_sig000004cd : STD_LOGIC; 
  signal blk00000003_sig000004cc : STD_LOGIC; 
  signal blk00000003_sig000004cb : STD_LOGIC; 
  signal blk00000003_sig000004ca : STD_LOGIC; 
  signal blk00000003_sig000004c9 : STD_LOGIC; 
  signal blk00000003_sig000004c8 : STD_LOGIC; 
  signal blk00000003_sig000004c7 : STD_LOGIC; 
  signal blk00000003_sig000004c6 : STD_LOGIC; 
  signal blk00000003_sig000004c5 : STD_LOGIC; 
  signal blk00000003_sig000004c4 : STD_LOGIC; 
  signal blk00000003_sig000004c3 : STD_LOGIC; 
  signal blk00000003_sig000004c2 : STD_LOGIC; 
  signal blk00000003_sig000004c1 : STD_LOGIC; 
  signal blk00000003_sig000004c0 : STD_LOGIC; 
  signal blk00000003_sig000004bf : STD_LOGIC; 
  signal blk00000003_sig000004be : STD_LOGIC; 
  signal blk00000003_sig000004bd : STD_LOGIC; 
  signal blk00000003_sig000004bc : STD_LOGIC; 
  signal blk00000003_sig000004bb : STD_LOGIC; 
  signal blk00000003_sig000004ba : STD_LOGIC; 
  signal blk00000003_sig000004b9 : STD_LOGIC; 
  signal blk00000003_sig000004b8 : STD_LOGIC; 
  signal blk00000003_sig000004b7 : STD_LOGIC; 
  signal blk00000003_sig000004b6 : STD_LOGIC; 
  signal blk00000003_sig000004b5 : STD_LOGIC; 
  signal blk00000003_sig000004b4 : STD_LOGIC; 
  signal blk00000003_sig000004b3 : STD_LOGIC; 
  signal blk00000003_sig000004b2 : STD_LOGIC; 
  signal blk00000003_sig000004b1 : STD_LOGIC; 
  signal blk00000003_sig000004b0 : STD_LOGIC; 
  signal blk00000003_sig000004af : STD_LOGIC; 
  signal blk00000003_sig000004ae : STD_LOGIC; 
  signal blk00000003_sig000004ad : STD_LOGIC; 
  signal blk00000003_sig000004ac : STD_LOGIC; 
  signal blk00000003_sig000004ab : STD_LOGIC; 
  signal blk00000003_sig000004aa : STD_LOGIC; 
  signal blk00000003_sig000004a9 : STD_LOGIC; 
  signal blk00000003_sig000004a8 : STD_LOGIC; 
  signal blk00000003_sig000004a7 : STD_LOGIC; 
  signal blk00000003_sig000004a6 : STD_LOGIC; 
  signal blk00000003_sig000004a5 : STD_LOGIC; 
  signal blk00000003_sig000004a4 : STD_LOGIC; 
  signal blk00000003_sig000004a3 : STD_LOGIC; 
  signal blk00000003_sig000004a2 : STD_LOGIC; 
  signal blk00000003_sig000004a1 : STD_LOGIC; 
  signal blk00000003_sig000004a0 : STD_LOGIC; 
  signal blk00000003_sig0000049f : STD_LOGIC; 
  signal blk00000003_sig0000049e : STD_LOGIC; 
  signal blk00000003_sig0000049d : STD_LOGIC; 
  signal blk00000003_sig0000049c : STD_LOGIC; 
  signal blk00000003_sig0000049b : STD_LOGIC; 
  signal blk00000003_sig0000049a : STD_LOGIC; 
  signal blk00000003_sig00000499 : STD_LOGIC; 
  signal blk00000003_sig00000498 : STD_LOGIC; 
  signal blk00000003_sig00000497 : STD_LOGIC; 
  signal blk00000003_sig00000496 : STD_LOGIC; 
  signal blk00000003_sig00000495 : STD_LOGIC; 
  signal blk00000003_sig00000494 : STD_LOGIC; 
  signal blk00000003_sig00000493 : STD_LOGIC; 
  signal blk00000003_sig00000492 : STD_LOGIC; 
  signal blk00000003_sig00000491 : STD_LOGIC; 
  signal blk00000003_sig00000490 : STD_LOGIC; 
  signal blk00000003_sig0000048f : STD_LOGIC; 
  signal blk00000003_sig0000048e : STD_LOGIC; 
  signal blk00000003_sig0000048d : STD_LOGIC; 
  signal blk00000003_sig0000048c : STD_LOGIC; 
  signal blk00000003_sig0000048b : STD_LOGIC; 
  signal blk00000003_sig0000048a : STD_LOGIC; 
  signal blk00000003_sig00000489 : STD_LOGIC; 
  signal blk00000003_sig00000488 : STD_LOGIC; 
  signal blk00000003_sig00000487 : STD_LOGIC; 
  signal blk00000003_sig00000486 : STD_LOGIC; 
  signal blk00000003_sig00000485 : STD_LOGIC; 
  signal blk00000003_sig00000484 : STD_LOGIC; 
  signal blk00000003_sig00000483 : STD_LOGIC; 
  signal blk00000003_sig00000482 : STD_LOGIC; 
  signal blk00000003_sig00000481 : STD_LOGIC; 
  signal blk00000003_sig00000480 : STD_LOGIC; 
  signal blk00000003_sig0000047f : STD_LOGIC; 
  signal blk00000003_sig0000047e : STD_LOGIC; 
  signal blk00000003_sig0000047d : STD_LOGIC; 
  signal blk00000003_sig0000047c : STD_LOGIC; 
  signal blk00000003_sig0000047b : STD_LOGIC; 
  signal blk00000003_sig0000047a : STD_LOGIC; 
  signal blk00000003_sig00000479 : STD_LOGIC; 
  signal blk00000003_sig00000478 : STD_LOGIC; 
  signal blk00000003_sig00000477 : STD_LOGIC; 
  signal blk00000003_sig00000476 : STD_LOGIC; 
  signal blk00000003_sig00000475 : STD_LOGIC; 
  signal blk00000003_sig00000474 : STD_LOGIC; 
  signal blk00000003_sig00000473 : STD_LOGIC; 
  signal blk00000003_sig00000472 : STD_LOGIC; 
  signal blk00000003_sig00000471 : STD_LOGIC; 
  signal blk00000003_sig00000470 : STD_LOGIC; 
  signal blk00000003_sig0000046f : STD_LOGIC; 
  signal blk00000003_sig0000046e : STD_LOGIC; 
  signal blk00000003_sig0000046d : STD_LOGIC; 
  signal blk00000003_sig0000046c : STD_LOGIC; 
  signal blk00000003_sig0000046b : STD_LOGIC; 
  signal blk00000003_sig0000046a : STD_LOGIC; 
  signal blk00000003_sig00000469 : STD_LOGIC; 
  signal blk00000003_sig00000468 : STD_LOGIC; 
  signal blk00000003_sig00000467 : STD_LOGIC; 
  signal blk00000003_sig00000466 : STD_LOGIC; 
  signal blk00000003_sig00000465 : STD_LOGIC; 
  signal blk00000003_sig00000464 : STD_LOGIC; 
  signal blk00000003_sig00000463 : STD_LOGIC; 
  signal blk00000003_sig00000462 : STD_LOGIC; 
  signal blk00000003_sig00000461 : STD_LOGIC; 
  signal blk00000003_sig00000460 : STD_LOGIC; 
  signal blk00000003_sig0000045f : STD_LOGIC; 
  signal blk00000003_sig0000045e : STD_LOGIC; 
  signal blk00000003_sig0000045d : STD_LOGIC; 
  signal blk00000003_sig0000045c : STD_LOGIC; 
  signal blk00000003_sig0000045b : STD_LOGIC; 
  signal blk00000003_sig0000045a : STD_LOGIC; 
  signal blk00000003_sig00000459 : STD_LOGIC; 
  signal blk00000003_sig00000458 : STD_LOGIC; 
  signal blk00000003_sig00000457 : STD_LOGIC; 
  signal blk00000003_sig00000456 : STD_LOGIC; 
  signal blk00000003_sig00000455 : STD_LOGIC; 
  signal blk00000003_sig00000454 : STD_LOGIC; 
  signal blk00000003_sig00000453 : STD_LOGIC; 
  signal blk00000003_sig00000452 : STD_LOGIC; 
  signal blk00000003_sig00000451 : STD_LOGIC; 
  signal blk00000003_sig00000450 : STD_LOGIC; 
  signal blk00000003_sig0000044f : STD_LOGIC; 
  signal blk00000003_sig0000044e : STD_LOGIC; 
  signal blk00000003_sig0000044d : STD_LOGIC; 
  signal blk00000003_sig0000044c : STD_LOGIC; 
  signal blk00000003_sig0000044b : STD_LOGIC; 
  signal blk00000003_sig0000044a : STD_LOGIC; 
  signal blk00000003_sig00000449 : STD_LOGIC; 
  signal blk00000003_sig00000448 : STD_LOGIC; 
  signal blk00000003_sig00000447 : STD_LOGIC; 
  signal blk00000003_sig00000446 : STD_LOGIC; 
  signal blk00000003_sig00000445 : STD_LOGIC; 
  signal blk00000003_sig00000444 : STD_LOGIC; 
  signal blk00000003_sig00000443 : STD_LOGIC; 
  signal blk00000003_sig00000442 : STD_LOGIC; 
  signal blk00000003_sig00000441 : STD_LOGIC; 
  signal blk00000003_sig00000440 : STD_LOGIC; 
  signal blk00000003_sig0000043f : STD_LOGIC; 
  signal blk00000003_sig0000043e : STD_LOGIC; 
  signal blk00000003_sig0000043d : STD_LOGIC; 
  signal blk00000003_sig0000043c : STD_LOGIC; 
  signal blk00000003_sig0000043b : STD_LOGIC; 
  signal blk00000003_sig0000043a : STD_LOGIC; 
  signal blk00000003_sig00000439 : STD_LOGIC; 
  signal blk00000003_sig00000438 : STD_LOGIC; 
  signal blk00000003_sig00000437 : STD_LOGIC; 
  signal blk00000003_sig00000436 : STD_LOGIC; 
  signal blk00000003_sig00000435 : STD_LOGIC; 
  signal blk00000003_sig00000434 : STD_LOGIC; 
  signal blk00000003_sig00000433 : STD_LOGIC; 
  signal blk00000003_sig00000432 : STD_LOGIC; 
  signal blk00000003_sig00000431 : STD_LOGIC; 
  signal blk00000003_sig00000430 : STD_LOGIC; 
  signal blk00000003_sig0000042f : STD_LOGIC; 
  signal blk00000003_sig0000042e : STD_LOGIC; 
  signal blk00000003_sig0000042d : STD_LOGIC; 
  signal blk00000003_sig0000042c : STD_LOGIC; 
  signal blk00000003_sig0000042b : STD_LOGIC; 
  signal blk00000003_sig0000042a : STD_LOGIC; 
  signal blk00000003_sig00000429 : STD_LOGIC; 
  signal blk00000003_sig00000428 : STD_LOGIC; 
  signal blk00000003_sig00000427 : STD_LOGIC; 
  signal blk00000003_sig00000426 : STD_LOGIC; 
  signal blk00000003_sig00000425 : STD_LOGIC; 
  signal blk00000003_sig00000424 : STD_LOGIC; 
  signal blk00000003_sig00000423 : STD_LOGIC; 
  signal blk00000003_sig00000422 : STD_LOGIC; 
  signal blk00000003_sig00000421 : STD_LOGIC; 
  signal blk00000003_sig00000420 : STD_LOGIC; 
  signal blk00000003_sig0000041f : STD_LOGIC; 
  signal blk00000003_sig0000041e : STD_LOGIC; 
  signal blk00000003_sig0000041d : STD_LOGIC; 
  signal blk00000003_sig0000041c : STD_LOGIC; 
  signal blk00000003_sig0000041b : STD_LOGIC; 
  signal blk00000003_sig0000041a : STD_LOGIC; 
  signal blk00000003_sig00000419 : STD_LOGIC; 
  signal blk00000003_sig00000418 : STD_LOGIC; 
  signal blk00000003_sig00000417 : STD_LOGIC; 
  signal blk00000003_sig00000416 : STD_LOGIC; 
  signal blk00000003_sig00000415 : STD_LOGIC; 
  signal blk00000003_sig00000414 : STD_LOGIC; 
  signal blk00000003_sig00000413 : STD_LOGIC; 
  signal blk00000003_sig00000412 : STD_LOGIC; 
  signal blk00000003_sig00000411 : STD_LOGIC; 
  signal blk00000003_sig00000410 : STD_LOGIC; 
  signal blk00000003_sig0000040f : STD_LOGIC; 
  signal blk00000003_sig0000040e : STD_LOGIC; 
  signal blk00000003_sig0000040d : STD_LOGIC; 
  signal blk00000003_sig0000040c : STD_LOGIC; 
  signal blk00000003_sig0000040b : STD_LOGIC; 
  signal blk00000003_sig0000040a : STD_LOGIC; 
  signal blk00000003_sig00000409 : STD_LOGIC; 
  signal blk00000003_sig00000408 : STD_LOGIC; 
  signal blk00000003_sig00000407 : STD_LOGIC; 
  signal blk00000003_sig00000406 : STD_LOGIC; 
  signal blk00000003_sig00000405 : STD_LOGIC; 
  signal blk00000003_sig00000404 : STD_LOGIC; 
  signal blk00000003_sig00000403 : STD_LOGIC; 
  signal blk00000003_sig00000402 : STD_LOGIC; 
  signal blk00000003_sig00000401 : STD_LOGIC; 
  signal blk00000003_sig00000400 : STD_LOGIC; 
  signal blk00000003_sig000003ff : STD_LOGIC; 
  signal blk00000003_sig000003fe : STD_LOGIC; 
  signal blk00000003_sig000003fd : STD_LOGIC; 
  signal blk00000003_sig000003fc : STD_LOGIC; 
  signal blk00000003_sig000003fb : STD_LOGIC; 
  signal blk00000003_sig000003fa : STD_LOGIC; 
  signal blk00000003_sig000003f9 : STD_LOGIC; 
  signal blk00000003_sig000003f8 : STD_LOGIC; 
  signal blk00000003_sig000003f7 : STD_LOGIC; 
  signal blk00000003_sig000003f6 : STD_LOGIC; 
  signal blk00000003_sig000003f5 : STD_LOGIC; 
  signal blk00000003_sig000003f4 : STD_LOGIC; 
  signal blk00000003_sig000003f3 : STD_LOGIC; 
  signal blk00000003_sig000003f2 : STD_LOGIC; 
  signal blk00000003_sig000003f1 : STD_LOGIC; 
  signal blk00000003_sig000003f0 : STD_LOGIC; 
  signal blk00000003_sig000003ef : STD_LOGIC; 
  signal blk00000003_sig000003ee : STD_LOGIC; 
  signal blk00000003_sig000003ed : STD_LOGIC; 
  signal blk00000003_sig000003ec : STD_LOGIC; 
  signal blk00000003_sig000003eb : STD_LOGIC; 
  signal blk00000003_sig000003ea : STD_LOGIC; 
  signal blk00000003_sig000003e9 : STD_LOGIC; 
  signal blk00000003_sig000003e8 : STD_LOGIC; 
  signal blk00000003_sig000003e7 : STD_LOGIC; 
  signal blk00000003_sig000003e6 : STD_LOGIC; 
  signal blk00000003_sig000003e5 : STD_LOGIC; 
  signal blk00000003_sig000003e4 : STD_LOGIC; 
  signal blk00000003_sig000003e3 : STD_LOGIC; 
  signal blk00000003_sig000003e2 : STD_LOGIC; 
  signal blk00000003_sig000003e1 : STD_LOGIC; 
  signal blk00000003_sig000003e0 : STD_LOGIC; 
  signal blk00000003_sig000003df : STD_LOGIC; 
  signal blk00000003_sig000003de : STD_LOGIC; 
  signal blk00000003_sig000003dd : STD_LOGIC; 
  signal blk00000003_sig000003dc : STD_LOGIC; 
  signal blk00000003_sig000003db : STD_LOGIC; 
  signal blk00000003_sig000003da : STD_LOGIC; 
  signal blk00000003_sig000003d9 : STD_LOGIC; 
  signal blk00000003_sig000003d8 : STD_LOGIC; 
  signal blk00000003_sig000003d7 : STD_LOGIC; 
  signal blk00000003_sig000003d6 : STD_LOGIC; 
  signal blk00000003_sig000003d5 : STD_LOGIC; 
  signal blk00000003_sig000003d4 : STD_LOGIC; 
  signal blk00000003_sig000003d3 : STD_LOGIC; 
  signal blk00000003_sig000003d2 : STD_LOGIC; 
  signal blk00000003_sig000003d1 : STD_LOGIC; 
  signal blk00000003_sig000003d0 : STD_LOGIC; 
  signal blk00000003_sig000003cf : STD_LOGIC; 
  signal blk00000003_sig000003ce : STD_LOGIC; 
  signal blk00000003_sig000003cd : STD_LOGIC; 
  signal blk00000003_sig000003cc : STD_LOGIC; 
  signal blk00000003_sig000003cb : STD_LOGIC; 
  signal blk00000003_sig000003ca : STD_LOGIC; 
  signal blk00000003_sig000003c9 : STD_LOGIC; 
  signal blk00000003_sig000003c8 : STD_LOGIC; 
  signal blk00000003_sig000003c7 : STD_LOGIC; 
  signal blk00000003_sig000003c6 : STD_LOGIC; 
  signal blk00000003_sig000003c5 : STD_LOGIC; 
  signal blk00000003_sig000003c4 : STD_LOGIC; 
  signal blk00000003_sig000003c3 : STD_LOGIC; 
  signal blk00000003_sig000003c2 : STD_LOGIC; 
  signal blk00000003_sig000003c1 : STD_LOGIC; 
  signal blk00000003_sig000003c0 : STD_LOGIC; 
  signal blk00000003_sig000003bf : STD_LOGIC; 
  signal blk00000003_sig000003be : STD_LOGIC; 
  signal blk00000003_sig000003bd : STD_LOGIC; 
  signal blk00000003_sig000003bc : STD_LOGIC; 
  signal blk00000003_sig000003bb : STD_LOGIC; 
  signal blk00000003_sig000003ba : STD_LOGIC; 
  signal blk00000003_sig000003b9 : STD_LOGIC; 
  signal blk00000003_sig000003b8 : STD_LOGIC; 
  signal blk00000003_sig000003b7 : STD_LOGIC; 
  signal blk00000003_sig000003b6 : STD_LOGIC; 
  signal blk00000003_sig000003b5 : STD_LOGIC; 
  signal blk00000003_sig000003b4 : STD_LOGIC; 
  signal blk00000003_sig000003b3 : STD_LOGIC; 
  signal blk00000003_sig000003b2 : STD_LOGIC; 
  signal blk00000003_sig000003b1 : STD_LOGIC; 
  signal blk00000003_sig000003b0 : STD_LOGIC; 
  signal blk00000003_sig000003af : STD_LOGIC; 
  signal blk00000003_sig000003ae : STD_LOGIC; 
  signal blk00000003_sig000003ad : STD_LOGIC; 
  signal blk00000003_sig000003ac : STD_LOGIC; 
  signal blk00000003_sig000003ab : STD_LOGIC; 
  signal blk00000003_sig000003aa : STD_LOGIC; 
  signal blk00000003_sig000003a9 : STD_LOGIC; 
  signal blk00000003_sig000003a8 : STD_LOGIC; 
  signal blk00000003_sig000003a7 : STD_LOGIC; 
  signal blk00000003_sig000003a6 : STD_LOGIC; 
  signal blk00000003_sig000003a5 : STD_LOGIC; 
  signal blk00000003_sig000003a4 : STD_LOGIC; 
  signal blk00000003_sig000003a3 : STD_LOGIC; 
  signal blk00000003_sig000003a2 : STD_LOGIC; 
  signal blk00000003_sig000003a1 : STD_LOGIC; 
  signal blk00000003_sig000003a0 : STD_LOGIC; 
  signal blk00000003_sig0000039f : STD_LOGIC; 
  signal blk00000003_sig0000039e : STD_LOGIC; 
  signal blk00000003_sig0000039d : STD_LOGIC; 
  signal blk00000003_sig0000039c : STD_LOGIC; 
  signal blk00000003_sig0000039b : STD_LOGIC; 
  signal blk00000003_sig0000039a : STD_LOGIC; 
  signal blk00000003_sig00000399 : STD_LOGIC; 
  signal blk00000003_sig00000398 : STD_LOGIC; 
  signal blk00000003_sig00000397 : STD_LOGIC; 
  signal blk00000003_sig00000396 : STD_LOGIC; 
  signal blk00000003_sig00000395 : STD_LOGIC; 
  signal blk00000003_sig00000394 : STD_LOGIC; 
  signal blk00000003_sig00000393 : STD_LOGIC; 
  signal blk00000003_sig00000392 : STD_LOGIC; 
  signal blk00000003_sig00000391 : STD_LOGIC; 
  signal blk00000003_sig00000390 : STD_LOGIC; 
  signal blk00000003_sig0000038f : STD_LOGIC; 
  signal blk00000003_sig0000038e : STD_LOGIC; 
  signal blk00000003_sig0000038d : STD_LOGIC; 
  signal blk00000003_sig0000038c : STD_LOGIC; 
  signal blk00000003_sig0000038b : STD_LOGIC; 
  signal blk00000003_sig0000038a : STD_LOGIC; 
  signal blk00000003_sig00000389 : STD_LOGIC; 
  signal blk00000003_sig00000388 : STD_LOGIC; 
  signal blk00000003_sig00000387 : STD_LOGIC; 
  signal blk00000003_sig00000386 : STD_LOGIC; 
  signal blk00000003_sig00000385 : STD_LOGIC; 
  signal blk00000003_sig00000384 : STD_LOGIC; 
  signal blk00000003_sig00000383 : STD_LOGIC; 
  signal blk00000003_sig00000382 : STD_LOGIC; 
  signal blk00000003_sig00000381 : STD_LOGIC; 
  signal blk00000003_sig00000380 : STD_LOGIC; 
  signal blk00000003_sig0000037f : STD_LOGIC; 
  signal blk00000003_sig0000037e : STD_LOGIC; 
  signal blk00000003_sig0000037d : STD_LOGIC; 
  signal blk00000003_sig0000037c : STD_LOGIC; 
  signal blk00000003_sig0000037b : STD_LOGIC; 
  signal blk00000003_sig0000037a : STD_LOGIC; 
  signal blk00000003_sig00000379 : STD_LOGIC; 
  signal blk00000003_sig00000378 : STD_LOGIC; 
  signal blk00000003_sig00000377 : STD_LOGIC; 
  signal blk00000003_sig00000376 : STD_LOGIC; 
  signal blk00000003_sig00000375 : STD_LOGIC; 
  signal blk00000003_sig00000374 : STD_LOGIC; 
  signal blk00000003_sig00000373 : STD_LOGIC; 
  signal blk00000003_sig00000372 : STD_LOGIC; 
  signal blk00000003_sig00000371 : STD_LOGIC; 
  signal blk00000003_sig00000370 : STD_LOGIC; 
  signal blk00000003_sig0000036f : STD_LOGIC; 
  signal blk00000003_sig0000036e : STD_LOGIC; 
  signal blk00000003_sig0000036d : STD_LOGIC; 
  signal blk00000003_sig0000036c : STD_LOGIC; 
  signal blk00000003_sig0000036b : STD_LOGIC; 
  signal blk00000003_sig0000036a : STD_LOGIC; 
  signal blk00000003_sig00000369 : STD_LOGIC; 
  signal blk00000003_sig00000368 : STD_LOGIC; 
  signal blk00000003_sig00000367 : STD_LOGIC; 
  signal blk00000003_sig00000366 : STD_LOGIC; 
  signal blk00000003_sig00000365 : STD_LOGIC; 
  signal blk00000003_sig00000364 : STD_LOGIC; 
  signal blk00000003_sig00000363 : STD_LOGIC; 
  signal blk00000003_sig00000362 : STD_LOGIC; 
  signal blk00000003_sig00000361 : STD_LOGIC; 
  signal blk00000003_sig00000360 : STD_LOGIC; 
  signal blk00000003_sig0000035f : STD_LOGIC; 
  signal blk00000003_sig0000035e : STD_LOGIC; 
  signal blk00000003_sig0000035d : STD_LOGIC; 
  signal blk00000003_sig0000035c : STD_LOGIC; 
  signal blk00000003_sig0000035b : STD_LOGIC; 
  signal blk00000003_sig0000035a : STD_LOGIC; 
  signal blk00000003_sig00000359 : STD_LOGIC; 
  signal blk00000003_sig00000358 : STD_LOGIC; 
  signal blk00000003_sig00000357 : STD_LOGIC; 
  signal blk00000003_sig00000356 : STD_LOGIC; 
  signal blk00000003_sig00000355 : STD_LOGIC; 
  signal blk00000003_sig00000354 : STD_LOGIC; 
  signal blk00000003_sig00000353 : STD_LOGIC; 
  signal blk00000003_sig00000352 : STD_LOGIC; 
  signal blk00000003_sig00000351 : STD_LOGIC; 
  signal blk00000003_sig00000350 : STD_LOGIC; 
  signal blk00000003_sig0000034f : STD_LOGIC; 
  signal blk00000003_sig0000034e : STD_LOGIC; 
  signal blk00000003_sig0000034d : STD_LOGIC; 
  signal blk00000003_sig0000034c : STD_LOGIC; 
  signal blk00000003_sig0000034b : STD_LOGIC; 
  signal blk00000003_sig0000034a : STD_LOGIC; 
  signal blk00000003_sig00000349 : STD_LOGIC; 
  signal blk00000003_sig00000348 : STD_LOGIC; 
  signal blk00000003_sig00000347 : STD_LOGIC; 
  signal blk00000003_sig00000346 : STD_LOGIC; 
  signal blk00000003_sig00000345 : STD_LOGIC; 
  signal blk00000003_sig00000344 : STD_LOGIC; 
  signal blk00000003_sig00000343 : STD_LOGIC; 
  signal blk00000003_sig00000342 : STD_LOGIC; 
  signal blk00000003_sig00000341 : STD_LOGIC; 
  signal blk00000003_sig00000340 : STD_LOGIC; 
  signal blk00000003_sig0000033f : STD_LOGIC; 
  signal blk00000003_sig0000033e : STD_LOGIC; 
  signal blk00000003_sig0000033d : STD_LOGIC; 
  signal blk00000003_sig0000033c : STD_LOGIC; 
  signal blk00000003_sig0000033b : STD_LOGIC; 
  signal blk00000003_sig0000033a : STD_LOGIC; 
  signal blk00000003_sig00000339 : STD_LOGIC; 
  signal blk00000003_sig00000338 : STD_LOGIC; 
  signal blk00000003_sig00000337 : STD_LOGIC; 
  signal blk00000003_sig00000336 : STD_LOGIC; 
  signal blk00000003_sig00000335 : STD_LOGIC; 
  signal blk00000003_sig00000334 : STD_LOGIC; 
  signal blk00000003_sig00000333 : STD_LOGIC; 
  signal blk00000003_sig00000332 : STD_LOGIC; 
  signal blk00000003_sig00000331 : STD_LOGIC; 
  signal blk00000003_sig00000330 : STD_LOGIC; 
  signal blk00000003_sig0000032f : STD_LOGIC; 
  signal blk00000003_sig0000032e : STD_LOGIC; 
  signal blk00000003_sig0000032d : STD_LOGIC; 
  signal blk00000003_sig0000032c : STD_LOGIC; 
  signal blk00000003_sig0000032b : STD_LOGIC; 
  signal blk00000003_sig0000032a : STD_LOGIC; 
  signal blk00000003_sig00000329 : STD_LOGIC; 
  signal blk00000003_sig00000328 : STD_LOGIC; 
  signal blk00000003_sig00000327 : STD_LOGIC; 
  signal blk00000003_sig00000326 : STD_LOGIC; 
  signal blk00000003_sig00000325 : STD_LOGIC; 
  signal blk00000003_sig00000324 : STD_LOGIC; 
  signal blk00000003_sig00000323 : STD_LOGIC; 
  signal blk00000003_sig00000322 : STD_LOGIC; 
  signal blk00000003_sig00000321 : STD_LOGIC; 
  signal blk00000003_sig00000320 : STD_LOGIC; 
  signal blk00000003_sig0000031f : STD_LOGIC; 
  signal blk00000003_sig0000031e : STD_LOGIC; 
  signal blk00000003_sig0000031d : STD_LOGIC; 
  signal blk00000003_sig0000031c : STD_LOGIC; 
  signal blk00000003_sig0000031b : STD_LOGIC; 
  signal blk00000003_sig0000031a : STD_LOGIC; 
  signal blk00000003_sig00000319 : STD_LOGIC; 
  signal blk00000003_sig00000318 : STD_LOGIC; 
  signal blk00000003_sig00000317 : STD_LOGIC; 
  signal blk00000003_sig00000316 : STD_LOGIC; 
  signal blk00000003_sig00000315 : STD_LOGIC; 
  signal blk00000003_sig00000314 : STD_LOGIC; 
  signal blk00000003_sig00000313 : STD_LOGIC; 
  signal blk00000003_sig00000312 : STD_LOGIC; 
  signal blk00000003_sig00000311 : STD_LOGIC; 
  signal blk00000003_sig00000310 : STD_LOGIC; 
  signal blk00000003_sig0000030f : STD_LOGIC; 
  signal blk00000003_sig0000030e : STD_LOGIC; 
  signal blk00000003_sig0000030d : STD_LOGIC; 
  signal blk00000003_sig0000030c : STD_LOGIC; 
  signal blk00000003_sig0000030b : STD_LOGIC; 
  signal blk00000003_sig0000030a : STD_LOGIC; 
  signal blk00000003_sig00000309 : STD_LOGIC; 
  signal blk00000003_sig00000308 : STD_LOGIC; 
  signal blk00000003_sig00000307 : STD_LOGIC; 
  signal blk00000003_sig00000306 : STD_LOGIC; 
  signal blk00000003_sig00000305 : STD_LOGIC; 
  signal blk00000003_sig00000304 : STD_LOGIC; 
  signal blk00000003_sig00000303 : STD_LOGIC; 
  signal blk00000003_sig00000302 : STD_LOGIC; 
  signal blk00000003_sig00000301 : STD_LOGIC; 
  signal blk00000003_sig00000300 : STD_LOGIC; 
  signal blk00000003_sig000002ff : STD_LOGIC; 
  signal blk00000003_sig000002fe : STD_LOGIC; 
  signal blk00000003_sig000002fd : STD_LOGIC; 
  signal blk00000003_sig000002fc : STD_LOGIC; 
  signal blk00000003_sig000002fb : STD_LOGIC; 
  signal blk00000003_sig000002fa : STD_LOGIC; 
  signal blk00000003_sig000002f9 : STD_LOGIC; 
  signal blk00000003_sig000002f8 : STD_LOGIC; 
  signal blk00000003_sig000002f7 : STD_LOGIC; 
  signal blk00000003_sig000002f6 : STD_LOGIC; 
  signal blk00000003_sig000002f5 : STD_LOGIC; 
  signal blk00000003_sig000002f4 : STD_LOGIC; 
  signal blk00000003_sig000002f3 : STD_LOGIC; 
  signal blk00000003_sig000002f2 : STD_LOGIC; 
  signal blk00000003_sig000002f1 : STD_LOGIC; 
  signal blk00000003_sig000002f0 : STD_LOGIC; 
  signal blk00000003_sig000002ef : STD_LOGIC; 
  signal blk00000003_sig000002ee : STD_LOGIC; 
  signal blk00000003_sig000002ed : STD_LOGIC; 
  signal blk00000003_sig000002ec : STD_LOGIC; 
  signal blk00000003_sig000002eb : STD_LOGIC; 
  signal blk00000003_sig000002ea : STD_LOGIC; 
  signal blk00000003_sig000002e9 : STD_LOGIC; 
  signal blk00000003_sig000002e8 : STD_LOGIC; 
  signal blk00000003_sig000002e7 : STD_LOGIC; 
  signal blk00000003_sig000002e6 : STD_LOGIC; 
  signal blk00000003_sig000002e5 : STD_LOGIC; 
  signal blk00000003_sig000002e4 : STD_LOGIC; 
  signal blk00000003_sig000002e3 : STD_LOGIC; 
  signal blk00000003_sig000002e2 : STD_LOGIC; 
  signal blk00000003_sig000002e1 : STD_LOGIC; 
  signal blk00000003_sig000002e0 : STD_LOGIC; 
  signal blk00000003_sig000002df : STD_LOGIC; 
  signal blk00000003_sig000002de : STD_LOGIC; 
  signal blk00000003_sig000002dd : STD_LOGIC; 
  signal blk00000003_sig000002dc : STD_LOGIC; 
  signal blk00000003_sig000002db : STD_LOGIC; 
  signal blk00000003_sig000002da : STD_LOGIC; 
  signal blk00000003_sig000002d9 : STD_LOGIC; 
  signal blk00000003_sig000002d8 : STD_LOGIC; 
  signal blk00000003_sig000002d7 : STD_LOGIC; 
  signal blk00000003_sig000002d6 : STD_LOGIC; 
  signal blk00000003_sig000002d5 : STD_LOGIC; 
  signal blk00000003_sig000002d4 : STD_LOGIC; 
  signal blk00000003_sig000002d3 : STD_LOGIC; 
  signal blk00000003_sig000002d2 : STD_LOGIC; 
  signal blk00000003_sig000002d1 : STD_LOGIC; 
  signal blk00000003_sig000002d0 : STD_LOGIC; 
  signal blk00000003_sig000002cf : STD_LOGIC; 
  signal blk00000003_sig000002ce : STD_LOGIC; 
  signal blk00000003_sig000002cd : STD_LOGIC; 
  signal blk00000003_sig000002cc : STD_LOGIC; 
  signal blk00000003_sig000002cb : STD_LOGIC; 
  signal blk00000003_sig000002ca : STD_LOGIC; 
  signal blk00000003_sig000002c9 : STD_LOGIC; 
  signal blk00000003_sig000002c8 : STD_LOGIC; 
  signal blk00000003_sig000002c7 : STD_LOGIC; 
  signal blk00000003_sig000002c6 : STD_LOGIC; 
  signal blk00000003_sig000002c5 : STD_LOGIC; 
  signal blk00000003_sig000002c4 : STD_LOGIC; 
  signal blk00000003_sig000002c3 : STD_LOGIC; 
  signal blk00000003_sig000002c2 : STD_LOGIC; 
  signal blk00000003_sig000002c1 : STD_LOGIC; 
  signal blk00000003_sig000002c0 : STD_LOGIC; 
  signal blk00000003_sig000002bf : STD_LOGIC; 
  signal blk00000003_sig000002be : STD_LOGIC; 
  signal blk00000003_sig000002bd : STD_LOGIC; 
  signal blk00000003_sig000002bc : STD_LOGIC; 
  signal blk00000003_sig000002bb : STD_LOGIC; 
  signal blk00000003_sig000002ba : STD_LOGIC; 
  signal blk00000003_sig000002b9 : STD_LOGIC; 
  signal blk00000003_sig000002b8 : STD_LOGIC; 
  signal blk00000003_sig000002b7 : STD_LOGIC; 
  signal blk00000003_sig000002b6 : STD_LOGIC; 
  signal blk00000003_sig000002b5 : STD_LOGIC; 
  signal blk00000003_sig000002b4 : STD_LOGIC; 
  signal blk00000003_sig000002b3 : STD_LOGIC; 
  signal blk00000003_sig000002b2 : STD_LOGIC; 
  signal blk00000003_sig000002b1 : STD_LOGIC; 
  signal blk00000003_sig000002b0 : STD_LOGIC; 
  signal blk00000003_sig000002af : STD_LOGIC; 
  signal blk00000003_sig000002ae : STD_LOGIC; 
  signal blk00000003_sig000002ad : STD_LOGIC; 
  signal blk00000003_sig000002ac : STD_LOGIC; 
  signal blk00000003_sig000002ab : STD_LOGIC; 
  signal blk00000003_sig000002aa : STD_LOGIC; 
  signal blk00000003_sig000002a9 : STD_LOGIC; 
  signal blk00000003_sig000002a8 : STD_LOGIC; 
  signal blk00000003_sig000002a7 : STD_LOGIC; 
  signal blk00000003_sig000002a6 : STD_LOGIC; 
  signal blk00000003_sig000002a5 : STD_LOGIC; 
  signal blk00000003_sig000002a4 : STD_LOGIC; 
  signal blk00000003_sig000002a3 : STD_LOGIC; 
  signal blk00000003_sig000002a2 : STD_LOGIC; 
  signal blk00000003_sig000002a1 : STD_LOGIC; 
  signal blk00000003_sig000002a0 : STD_LOGIC; 
  signal blk00000003_sig0000029f : STD_LOGIC; 
  signal blk00000003_sig0000029e : STD_LOGIC; 
  signal blk00000003_sig0000029d : STD_LOGIC; 
  signal blk00000003_sig0000029c : STD_LOGIC; 
  signal blk00000003_sig0000029b : STD_LOGIC; 
  signal blk00000003_sig0000029a : STD_LOGIC; 
  signal blk00000003_sig00000299 : STD_LOGIC; 
  signal blk00000003_sig00000298 : STD_LOGIC; 
  signal blk00000003_sig00000297 : STD_LOGIC; 
  signal blk00000003_sig00000296 : STD_LOGIC; 
  signal blk00000003_sig00000295 : STD_LOGIC; 
  signal blk00000003_sig00000294 : STD_LOGIC; 
  signal blk00000003_sig00000293 : STD_LOGIC; 
  signal blk00000003_sig00000292 : STD_LOGIC; 
  signal blk00000003_sig00000291 : STD_LOGIC; 
  signal blk00000003_sig00000290 : STD_LOGIC; 
  signal blk00000003_sig0000028f : STD_LOGIC; 
  signal blk00000003_sig0000028e : STD_LOGIC; 
  signal blk00000003_sig0000028d : STD_LOGIC; 
  signal blk00000003_sig0000028c : STD_LOGIC; 
  signal blk00000003_sig0000028b : STD_LOGIC; 
  signal blk00000003_sig0000028a : STD_LOGIC; 
  signal blk00000003_sig00000289 : STD_LOGIC; 
  signal blk00000003_sig00000288 : STD_LOGIC; 
  signal blk00000003_sig00000287 : STD_LOGIC; 
  signal blk00000003_sig00000286 : STD_LOGIC; 
  signal blk00000003_sig00000285 : STD_LOGIC; 
  signal blk00000003_sig00000284 : STD_LOGIC; 
  signal blk00000003_sig00000283 : STD_LOGIC; 
  signal blk00000003_sig00000282 : STD_LOGIC; 
  signal blk00000003_sig00000281 : STD_LOGIC; 
  signal blk00000003_sig00000280 : STD_LOGIC; 
  signal blk00000003_sig0000027f : STD_LOGIC; 
  signal blk00000003_sig0000027e : STD_LOGIC; 
  signal blk00000003_sig0000027d : STD_LOGIC; 
  signal blk00000003_sig0000027c : STD_LOGIC; 
  signal blk00000003_sig0000027b : STD_LOGIC; 
  signal blk00000003_sig0000027a : STD_LOGIC; 
  signal blk00000003_sig00000279 : STD_LOGIC; 
  signal blk00000003_sig00000278 : STD_LOGIC; 
  signal blk00000003_sig00000277 : STD_LOGIC; 
  signal blk00000003_sig00000276 : STD_LOGIC; 
  signal blk00000003_sig00000275 : STD_LOGIC; 
  signal blk00000003_sig00000274 : STD_LOGIC; 
  signal blk00000003_sig00000273 : STD_LOGIC; 
  signal blk00000003_sig00000272 : STD_LOGIC; 
  signal blk00000003_sig00000271 : STD_LOGIC; 
  signal blk00000003_sig00000270 : STD_LOGIC; 
  signal blk00000003_sig0000026f : STD_LOGIC; 
  signal blk00000003_sig0000026e : STD_LOGIC; 
  signal blk00000003_sig0000026d : STD_LOGIC; 
  signal blk00000003_sig0000026c : STD_LOGIC; 
  signal blk00000003_sig0000026b : STD_LOGIC; 
  signal blk00000003_sig0000026a : STD_LOGIC; 
  signal blk00000003_sig00000269 : STD_LOGIC; 
  signal blk00000003_sig00000268 : STD_LOGIC; 
  signal blk00000003_sig00000267 : STD_LOGIC; 
  signal blk00000003_sig00000266 : STD_LOGIC; 
  signal blk00000003_sig00000265 : STD_LOGIC; 
  signal blk00000003_sig00000264 : STD_LOGIC; 
  signal blk00000003_sig00000263 : STD_LOGIC; 
  signal blk00000003_sig00000262 : STD_LOGIC; 
  signal blk00000003_sig00000261 : STD_LOGIC; 
  signal blk00000003_sig00000260 : STD_LOGIC; 
  signal blk00000003_sig0000025f : STD_LOGIC; 
  signal blk00000003_sig0000025e : STD_LOGIC; 
  signal blk00000003_sig0000025d : STD_LOGIC; 
  signal blk00000003_sig0000025c : STD_LOGIC; 
  signal blk00000003_sig0000025b : STD_LOGIC; 
  signal blk00000003_sig0000025a : STD_LOGIC; 
  signal blk00000003_sig00000259 : STD_LOGIC; 
  signal blk00000003_sig00000258 : STD_LOGIC; 
  signal blk00000003_sig00000257 : STD_LOGIC; 
  signal blk00000003_sig00000256 : STD_LOGIC; 
  signal blk00000003_sig00000255 : STD_LOGIC; 
  signal blk00000003_sig00000254 : STD_LOGIC; 
  signal blk00000003_sig00000253 : STD_LOGIC; 
  signal blk00000003_sig00000252 : STD_LOGIC; 
  signal blk00000003_sig00000251 : STD_LOGIC; 
  signal blk00000003_sig00000250 : STD_LOGIC; 
  signal blk00000003_sig0000024f : STD_LOGIC; 
  signal blk00000003_sig0000024e : STD_LOGIC; 
  signal blk00000003_sig0000024d : STD_LOGIC; 
  signal blk00000003_sig0000024c : STD_LOGIC; 
  signal blk00000003_sig0000024b : STD_LOGIC; 
  signal blk00000003_sig0000024a : STD_LOGIC; 
  signal blk00000003_sig00000249 : STD_LOGIC; 
  signal blk00000003_sig00000248 : STD_LOGIC; 
  signal blk00000003_sig00000247 : STD_LOGIC; 
  signal blk00000003_sig00000246 : STD_LOGIC; 
  signal blk00000003_sig00000245 : STD_LOGIC; 
  signal blk00000003_sig00000244 : STD_LOGIC; 
  signal blk00000003_sig00000243 : STD_LOGIC; 
  signal blk00000003_sig00000242 : STD_LOGIC; 
  signal blk00000003_sig00000241 : STD_LOGIC; 
  signal blk00000003_sig00000240 : STD_LOGIC; 
  signal blk00000003_sig0000023f : STD_LOGIC; 
  signal blk00000003_sig0000023e : STD_LOGIC; 
  signal blk00000003_sig0000023d : STD_LOGIC; 
  signal blk00000003_sig0000023c : STD_LOGIC; 
  signal blk00000003_sig0000023b : STD_LOGIC; 
  signal blk00000003_sig0000023a : STD_LOGIC; 
  signal blk00000003_sig00000239 : STD_LOGIC; 
  signal blk00000003_sig00000238 : STD_LOGIC; 
  signal blk00000003_sig00000237 : STD_LOGIC; 
  signal blk00000003_sig00000236 : STD_LOGIC; 
  signal blk00000003_sig00000235 : STD_LOGIC; 
  signal blk00000003_sig00000234 : STD_LOGIC; 
  signal blk00000003_sig00000233 : STD_LOGIC; 
  signal blk00000003_sig00000232 : STD_LOGIC; 
  signal blk00000003_sig00000231 : STD_LOGIC; 
  signal blk00000003_sig00000230 : STD_LOGIC; 
  signal blk00000003_sig0000022f : STD_LOGIC; 
  signal blk00000003_sig0000022e : STD_LOGIC; 
  signal blk00000003_sig0000022d : STD_LOGIC; 
  signal blk00000003_sig0000022c : STD_LOGIC; 
  signal blk00000003_sig0000022b : STD_LOGIC; 
  signal blk00000003_sig0000022a : STD_LOGIC; 
  signal blk00000003_sig00000229 : STD_LOGIC; 
  signal blk00000003_sig00000228 : STD_LOGIC; 
  signal blk00000003_sig00000227 : STD_LOGIC; 
  signal blk00000003_sig00000226 : STD_LOGIC; 
  signal blk00000003_sig00000225 : STD_LOGIC; 
  signal blk00000003_sig00000224 : STD_LOGIC; 
  signal blk00000003_sig00000223 : STD_LOGIC; 
  signal blk00000003_sig00000222 : STD_LOGIC; 
  signal blk00000003_sig00000221 : STD_LOGIC; 
  signal blk00000003_sig00000220 : STD_LOGIC; 
  signal blk00000003_sig0000021f : STD_LOGIC; 
  signal blk00000003_sig0000021e : STD_LOGIC; 
  signal blk00000003_sig0000021d : STD_LOGIC; 
  signal blk00000003_sig0000021c : STD_LOGIC; 
  signal blk00000003_sig0000021b : STD_LOGIC; 
  signal blk00000003_sig0000021a : STD_LOGIC; 
  signal blk00000003_sig00000219 : STD_LOGIC; 
  signal blk00000003_sig00000218 : STD_LOGIC; 
  signal blk00000003_sig00000217 : STD_LOGIC; 
  signal blk00000003_sig00000216 : STD_LOGIC; 
  signal blk00000003_sig00000215 : STD_LOGIC; 
  signal blk00000003_sig00000214 : STD_LOGIC; 
  signal blk00000003_sig00000213 : STD_LOGIC; 
  signal blk00000003_sig00000212 : STD_LOGIC; 
  signal blk00000003_sig00000211 : STD_LOGIC; 
  signal blk00000003_sig00000210 : STD_LOGIC; 
  signal blk00000003_sig0000020f : STD_LOGIC; 
  signal blk00000003_sig0000020e : STD_LOGIC; 
  signal blk00000003_sig0000020d : STD_LOGIC; 
  signal blk00000003_sig0000020c : STD_LOGIC; 
  signal blk00000003_sig0000020b : STD_LOGIC; 
  signal blk00000003_sig0000020a : STD_LOGIC; 
  signal blk00000003_sig00000209 : STD_LOGIC; 
  signal blk00000003_sig00000208 : STD_LOGIC; 
  signal blk00000003_sig00000207 : STD_LOGIC; 
  signal blk00000003_sig00000206 : STD_LOGIC; 
  signal blk00000003_sig00000205 : STD_LOGIC; 
  signal blk00000003_sig00000204 : STD_LOGIC; 
  signal blk00000003_sig00000203 : STD_LOGIC; 
  signal blk00000003_sig00000202 : STD_LOGIC; 
  signal blk00000003_sig00000201 : STD_LOGIC; 
  signal blk00000003_sig00000200 : STD_LOGIC; 
  signal blk00000003_sig000001ff : STD_LOGIC; 
  signal blk00000003_sig000001fe : STD_LOGIC; 
  signal blk00000003_sig000001fd : STD_LOGIC; 
  signal blk00000003_sig000001fc : STD_LOGIC; 
  signal blk00000003_sig000001fb : STD_LOGIC; 
  signal blk00000003_sig000001fa : STD_LOGIC; 
  signal blk00000003_sig000001f9 : STD_LOGIC; 
  signal blk00000003_sig000001f8 : STD_LOGIC; 
  signal blk00000003_sig000001f7 : STD_LOGIC; 
  signal blk00000003_sig000001f6 : STD_LOGIC; 
  signal blk00000003_sig000001f5 : STD_LOGIC; 
  signal blk00000003_sig000001f4 : STD_LOGIC; 
  signal blk00000003_sig000001f3 : STD_LOGIC; 
  signal blk00000003_sig000001f2 : STD_LOGIC; 
  signal blk00000003_sig000001f1 : STD_LOGIC; 
  signal blk00000003_sig000001f0 : STD_LOGIC; 
  signal blk00000003_sig000001ef : STD_LOGIC; 
  signal blk00000003_sig000001ee : STD_LOGIC; 
  signal blk00000003_sig000001ed : STD_LOGIC; 
  signal blk00000003_sig000001ec : STD_LOGIC; 
  signal blk00000003_sig000001eb : STD_LOGIC; 
  signal blk00000003_sig000001ea : STD_LOGIC; 
  signal blk00000003_sig000001e9 : STD_LOGIC; 
  signal blk00000003_sig000001e8 : STD_LOGIC; 
  signal blk00000003_sig000001e7 : STD_LOGIC; 
  signal blk00000003_sig000001e6 : STD_LOGIC; 
  signal blk00000003_sig000001e5 : STD_LOGIC; 
  signal blk00000003_sig000001e4 : STD_LOGIC; 
  signal blk00000003_sig000001e3 : STD_LOGIC; 
  signal blk00000003_sig000001e2 : STD_LOGIC; 
  signal blk00000003_sig000001e1 : STD_LOGIC; 
  signal blk00000003_sig000001e0 : STD_LOGIC; 
  signal blk00000003_sig000001df : STD_LOGIC; 
  signal blk00000003_sig000001de : STD_LOGIC; 
  signal blk00000003_sig000001dd : STD_LOGIC; 
  signal blk00000003_sig000001dc : STD_LOGIC; 
  signal blk00000003_sig000001db : STD_LOGIC; 
  signal blk00000003_sig000001da : STD_LOGIC; 
  signal blk00000003_sig000001d9 : STD_LOGIC; 
  signal blk00000003_sig000001d8 : STD_LOGIC; 
  signal blk00000003_sig000001d7 : STD_LOGIC; 
  signal blk00000003_sig000001d6 : STD_LOGIC; 
  signal blk00000003_sig000001d5 : STD_LOGIC; 
  signal blk00000003_sig000001d4 : STD_LOGIC; 
  signal blk00000003_sig000001d3 : STD_LOGIC; 
  signal blk00000003_sig000001d2 : STD_LOGIC; 
  signal blk00000003_sig000001d1 : STD_LOGIC; 
  signal blk00000003_sig000001d0 : STD_LOGIC; 
  signal blk00000003_sig000001cf : STD_LOGIC; 
  signal blk00000003_sig000001ce : STD_LOGIC; 
  signal blk00000003_sig000001cd : STD_LOGIC; 
  signal blk00000003_sig000001cc : STD_LOGIC; 
  signal blk00000003_sig000001cb : STD_LOGIC; 
  signal blk00000003_sig000001ca : STD_LOGIC; 
  signal blk00000003_sig000001c9 : STD_LOGIC; 
  signal blk00000003_sig000001c8 : STD_LOGIC; 
  signal blk00000003_sig000001c7 : STD_LOGIC; 
  signal blk00000003_sig000001c6 : STD_LOGIC; 
  signal blk00000003_sig000001c5 : STD_LOGIC; 
  signal blk00000003_sig000001c4 : STD_LOGIC; 
  signal blk00000003_sig000001c3 : STD_LOGIC; 
  signal blk00000003_sig000001c2 : STD_LOGIC; 
  signal blk00000003_sig000001c1 : STD_LOGIC; 
  signal blk00000003_sig000001c0 : STD_LOGIC; 
  signal blk00000003_sig000001bf : STD_LOGIC; 
  signal blk00000003_sig000001be : STD_LOGIC; 
  signal blk00000003_sig000001bd : STD_LOGIC; 
  signal blk00000003_sig000001bc : STD_LOGIC; 
  signal blk00000003_sig000001bb : STD_LOGIC; 
  signal blk00000003_sig000001ba : STD_LOGIC; 
  signal blk00000003_sig000001b9 : STD_LOGIC; 
  signal blk00000003_sig000001b8 : STD_LOGIC; 
  signal blk00000003_sig000001b7 : STD_LOGIC; 
  signal blk00000003_sig000001b6 : STD_LOGIC; 
  signal blk00000003_sig000001b5 : STD_LOGIC; 
  signal blk00000003_sig000001b4 : STD_LOGIC; 
  signal blk00000003_sig000001b3 : STD_LOGIC; 
  signal blk00000003_sig000001b2 : STD_LOGIC; 
  signal blk00000003_sig000001b1 : STD_LOGIC; 
  signal blk00000003_sig000001b0 : STD_LOGIC; 
  signal blk00000003_sig000001af : STD_LOGIC; 
  signal blk00000003_sig000001ae : STD_LOGIC; 
  signal blk00000003_sig000001ad : STD_LOGIC; 
  signal blk00000003_sig000001ac : STD_LOGIC; 
  signal blk00000003_sig000001ab : STD_LOGIC; 
  signal blk00000003_sig000001aa : STD_LOGIC; 
  signal blk00000003_sig000001a9 : STD_LOGIC; 
  signal blk00000003_sig000001a8 : STD_LOGIC; 
  signal blk00000003_sig000001a7 : STD_LOGIC; 
  signal blk00000003_sig000001a6 : STD_LOGIC; 
  signal blk00000003_sig000001a5 : STD_LOGIC; 
  signal blk00000003_sig000001a4 : STD_LOGIC; 
  signal blk00000003_sig000001a3 : STD_LOGIC; 
  signal blk00000003_sig000001a2 : STD_LOGIC; 
  signal blk00000003_sig000001a1 : STD_LOGIC; 
  signal blk00000003_sig000001a0 : STD_LOGIC; 
  signal blk00000003_sig0000019f : STD_LOGIC; 
  signal blk00000003_sig0000019e : STD_LOGIC; 
  signal blk00000003_sig0000019d : STD_LOGIC; 
  signal blk00000003_sig0000019c : STD_LOGIC; 
  signal blk00000003_sig0000019b : STD_LOGIC; 
  signal blk00000003_sig0000019a : STD_LOGIC; 
  signal blk00000003_sig00000199 : STD_LOGIC; 
  signal blk00000003_sig00000198 : STD_LOGIC; 
  signal blk00000003_sig00000197 : STD_LOGIC; 
  signal blk00000003_sig00000196 : STD_LOGIC; 
  signal blk00000003_sig00000195 : STD_LOGIC; 
  signal blk00000003_sig00000194 : STD_LOGIC; 
  signal blk00000003_sig00000193 : STD_LOGIC; 
  signal blk00000003_sig00000192 : STD_LOGIC; 
  signal blk00000003_sig00000191 : STD_LOGIC; 
  signal blk00000003_sig00000190 : STD_LOGIC; 
  signal blk00000003_sig0000018f : STD_LOGIC; 
  signal blk00000003_sig0000018e : STD_LOGIC; 
  signal blk00000003_sig0000018d : STD_LOGIC; 
  signal blk00000003_sig0000018c : STD_LOGIC; 
  signal blk00000003_sig0000018b : STD_LOGIC; 
  signal blk00000003_sig0000018a : STD_LOGIC; 
  signal blk00000003_sig00000189 : STD_LOGIC; 
  signal blk00000003_sig00000188 : STD_LOGIC; 
  signal blk00000003_sig00000187 : STD_LOGIC; 
  signal blk00000003_sig00000186 : STD_LOGIC; 
  signal blk00000003_sig00000185 : STD_LOGIC; 
  signal blk00000003_sig00000184 : STD_LOGIC; 
  signal blk00000003_sig00000183 : STD_LOGIC; 
  signal blk00000003_sig00000182 : STD_LOGIC; 
  signal blk00000003_sig00000181 : STD_LOGIC; 
  signal blk00000003_sig00000180 : STD_LOGIC; 
  signal blk00000003_sig0000017f : STD_LOGIC; 
  signal blk00000003_sig0000017e : STD_LOGIC; 
  signal blk00000003_sig0000017d : STD_LOGIC; 
  signal blk00000003_sig0000017c : STD_LOGIC; 
  signal blk00000003_sig0000017b : STD_LOGIC; 
  signal blk00000003_sig0000017a : STD_LOGIC; 
  signal blk00000003_sig00000179 : STD_LOGIC; 
  signal blk00000003_sig00000178 : STD_LOGIC; 
  signal blk00000003_sig00000177 : STD_LOGIC; 
  signal blk00000003_sig00000176 : STD_LOGIC; 
  signal blk00000003_sig00000175 : STD_LOGIC; 
  signal blk00000003_sig00000174 : STD_LOGIC; 
  signal blk00000003_sig00000173 : STD_LOGIC; 
  signal blk00000003_sig00000172 : STD_LOGIC; 
  signal blk00000003_sig00000171 : STD_LOGIC; 
  signal blk00000003_sig00000170 : STD_LOGIC; 
  signal blk00000003_sig0000016f : STD_LOGIC; 
  signal blk00000003_sig0000016e : STD_LOGIC; 
  signal blk00000003_sig0000016d : STD_LOGIC; 
  signal blk00000003_sig0000016c : STD_LOGIC; 
  signal blk00000003_sig0000016b : STD_LOGIC; 
  signal blk00000003_sig0000016a : STD_LOGIC; 
  signal blk00000003_sig00000169 : STD_LOGIC; 
  signal blk00000003_sig00000168 : STD_LOGIC; 
  signal blk00000003_sig00000167 : STD_LOGIC; 
  signal blk00000003_sig00000166 : STD_LOGIC; 
  signal blk00000003_sig00000165 : STD_LOGIC; 
  signal blk00000003_sig00000164 : STD_LOGIC; 
  signal blk00000003_sig00000163 : STD_LOGIC; 
  signal blk00000003_sig00000162 : STD_LOGIC; 
  signal blk00000003_sig00000161 : STD_LOGIC; 
  signal blk00000003_sig00000160 : STD_LOGIC; 
  signal blk00000003_sig0000015f : STD_LOGIC; 
  signal blk00000003_sig0000015e : STD_LOGIC; 
  signal blk00000003_sig0000015d : STD_LOGIC; 
  signal blk00000003_sig0000015c : STD_LOGIC; 
  signal blk00000003_sig0000015b : STD_LOGIC; 
  signal blk00000003_sig0000015a : STD_LOGIC; 
  signal blk00000003_sig00000159 : STD_LOGIC; 
  signal blk00000003_sig00000158 : STD_LOGIC; 
  signal blk00000003_sig00000157 : STD_LOGIC; 
  signal blk00000003_sig00000156 : STD_LOGIC; 
  signal blk00000003_sig00000155 : STD_LOGIC; 
  signal blk00000003_sig00000154 : STD_LOGIC; 
  signal blk00000003_sig00000153 : STD_LOGIC; 
  signal blk00000003_sig00000152 : STD_LOGIC; 
  signal blk00000003_sig00000151 : STD_LOGIC; 
  signal blk00000003_sig00000150 : STD_LOGIC; 
  signal blk00000003_sig0000014f : STD_LOGIC; 
  signal blk00000003_sig0000014e : STD_LOGIC; 
  signal blk00000003_sig0000014d : STD_LOGIC; 
  signal blk00000003_sig0000014c : STD_LOGIC; 
  signal blk00000003_sig0000014b : STD_LOGIC; 
  signal blk00000003_sig0000014a : STD_LOGIC; 
  signal blk00000003_sig00000149 : STD_LOGIC; 
  signal blk00000003_sig00000148 : STD_LOGIC; 
  signal blk00000003_sig00000147 : STD_LOGIC; 
  signal blk00000003_sig00000146 : STD_LOGIC; 
  signal blk00000003_sig00000145 : STD_LOGIC; 
  signal blk00000003_sig00000144 : STD_LOGIC; 
  signal blk00000003_sig00000143 : STD_LOGIC; 
  signal blk00000003_sig00000142 : STD_LOGIC; 
  signal blk00000003_sig00000141 : STD_LOGIC; 
  signal blk00000003_sig00000140 : STD_LOGIC; 
  signal blk00000003_sig0000013f : STD_LOGIC; 
  signal blk00000003_sig0000013e : STD_LOGIC; 
  signal blk00000003_sig0000013d : STD_LOGIC; 
  signal blk00000003_sig0000013c : STD_LOGIC; 
  signal blk00000003_sig0000013b : STD_LOGIC; 
  signal blk00000003_sig0000013a : STD_LOGIC; 
  signal blk00000003_sig00000139 : STD_LOGIC; 
  signal blk00000003_sig00000138 : STD_LOGIC; 
  signal blk00000003_sig00000137 : STD_LOGIC; 
  signal blk00000003_sig00000136 : STD_LOGIC; 
  signal blk00000003_sig00000135 : STD_LOGIC; 
  signal blk00000003_sig00000134 : STD_LOGIC; 
  signal blk00000003_sig00000133 : STD_LOGIC; 
  signal blk00000003_sig00000132 : STD_LOGIC; 
  signal blk00000003_sig00000131 : STD_LOGIC; 
  signal blk00000003_sig00000130 : STD_LOGIC; 
  signal blk00000003_sig0000012f : STD_LOGIC; 
  signal blk00000003_sig0000012e : STD_LOGIC; 
  signal blk00000003_sig0000012d : STD_LOGIC; 
  signal blk00000003_sig0000012c : STD_LOGIC; 
  signal blk00000003_sig0000012b : STD_LOGIC; 
  signal blk00000003_sig0000012a : STD_LOGIC; 
  signal blk00000003_sig00000129 : STD_LOGIC; 
  signal blk00000003_sig00000128 : STD_LOGIC; 
  signal blk00000003_sig00000127 : STD_LOGIC; 
  signal blk00000003_sig00000126 : STD_LOGIC; 
  signal blk00000003_sig00000125 : STD_LOGIC; 
  signal blk00000003_sig00000124 : STD_LOGIC; 
  signal blk00000003_sig00000123 : STD_LOGIC; 
  signal blk00000003_sig00000122 : STD_LOGIC; 
  signal blk00000003_sig00000121 : STD_LOGIC; 
  signal blk00000003_sig00000120 : STD_LOGIC; 
  signal blk00000003_sig0000011f : STD_LOGIC; 
  signal blk00000003_sig0000011e : STD_LOGIC; 
  signal blk00000003_sig0000011d : STD_LOGIC; 
  signal blk00000003_sig0000011c : STD_LOGIC; 
  signal blk00000003_sig0000011b : STD_LOGIC; 
  signal blk00000003_sig0000011a : STD_LOGIC; 
  signal blk00000003_sig00000119 : STD_LOGIC; 
  signal blk00000003_sig00000118 : STD_LOGIC; 
  signal blk00000003_sig00000117 : STD_LOGIC; 
  signal blk00000003_sig00000116 : STD_LOGIC; 
  signal blk00000003_sig00000115 : STD_LOGIC; 
  signal blk00000003_sig00000114 : STD_LOGIC; 
  signal blk00000003_sig00000113 : STD_LOGIC; 
  signal blk00000003_sig00000112 : STD_LOGIC; 
  signal blk00000003_sig00000111 : STD_LOGIC; 
  signal blk00000003_sig00000110 : STD_LOGIC; 
  signal blk00000003_sig0000010f : STD_LOGIC; 
  signal blk00000003_sig0000010e : STD_LOGIC; 
  signal blk00000003_sig0000010d : STD_LOGIC; 
  signal blk00000003_sig0000010c : STD_LOGIC; 
  signal blk00000003_sig0000010b : STD_LOGIC; 
  signal blk00000003_sig0000010a : STD_LOGIC; 
  signal blk00000003_sig00000109 : STD_LOGIC; 
  signal blk00000003_sig00000108 : STD_LOGIC; 
  signal blk00000003_sig00000107 : STD_LOGIC; 
  signal blk00000003_sig00000106 : STD_LOGIC; 
  signal blk00000003_sig00000105 : STD_LOGIC; 
  signal blk00000003_sig00000104 : STD_LOGIC; 
  signal blk00000003_sig00000103 : STD_LOGIC; 
  signal blk00000003_sig00000102 : STD_LOGIC; 
  signal blk00000003_sig00000101 : STD_LOGIC; 
  signal blk00000003_sig00000100 : STD_LOGIC; 
  signal blk00000003_sig000000ff : STD_LOGIC; 
  signal blk00000003_sig000000fe : STD_LOGIC; 
  signal blk00000003_sig000000fd : STD_LOGIC; 
  signal blk00000003_sig000000fc : STD_LOGIC; 
  signal blk00000003_sig000000fb : STD_LOGIC; 
  signal blk00000003_sig000000fa : STD_LOGIC; 
  signal blk00000003_sig000000f9 : STD_LOGIC; 
  signal blk00000003_sig000000f8 : STD_LOGIC; 
  signal blk00000003_sig000000f7 : STD_LOGIC; 
  signal blk00000003_sig000000f6 : STD_LOGIC; 
  signal blk00000003_sig000000f5 : STD_LOGIC; 
  signal blk00000003_sig000000f4 : STD_LOGIC; 
  signal blk00000003_sig000000f3 : STD_LOGIC; 
  signal blk00000003_sig000000f2 : STD_LOGIC; 
  signal blk00000003_sig000000f1 : STD_LOGIC; 
  signal blk00000003_sig000000f0 : STD_LOGIC; 
  signal blk00000003_sig000000ef : STD_LOGIC; 
  signal blk00000003_sig000000ee : STD_LOGIC; 
  signal blk00000003_sig000000ed : STD_LOGIC; 
  signal blk00000003_sig000000ec : STD_LOGIC; 
  signal blk00000003_sig000000eb : STD_LOGIC; 
  signal blk00000003_sig000000ea : STD_LOGIC; 
  signal blk00000003_sig000000e9 : STD_LOGIC; 
  signal blk00000003_sig000000e8 : STD_LOGIC; 
  signal blk00000003_sig000000e7 : STD_LOGIC; 
  signal blk00000003_sig000000e6 : STD_LOGIC; 
  signal blk00000003_sig000000e5 : STD_LOGIC; 
  signal blk00000003_sig000000e4 : STD_LOGIC; 
  signal blk00000003_sig000000e3 : STD_LOGIC; 
  signal blk00000003_sig000000e2 : STD_LOGIC; 
  signal blk00000003_sig000000e1 : STD_LOGIC; 
  signal blk00000003_sig000000e0 : STD_LOGIC; 
  signal blk00000003_sig000000df : STD_LOGIC; 
  signal blk00000003_sig000000de : STD_LOGIC; 
  signal blk00000003_sig000000dd : STD_LOGIC; 
  signal blk00000003_sig000000dc : STD_LOGIC; 
  signal blk00000003_sig000000db : STD_LOGIC; 
  signal blk00000003_sig000000da : STD_LOGIC; 
  signal blk00000003_sig000000d9 : STD_LOGIC; 
  signal blk00000003_sig000000d8 : STD_LOGIC; 
  signal blk00000003_sig000000d7 : STD_LOGIC; 
  signal blk00000003_sig000000d6 : STD_LOGIC; 
  signal blk00000003_sig000000d5 : STD_LOGIC; 
  signal blk00000003_sig000000d4 : STD_LOGIC; 
  signal blk00000003_sig000000d3 : STD_LOGIC; 
  signal blk00000003_sig000000d2 : STD_LOGIC; 
  signal blk00000003_sig000000d1 : STD_LOGIC; 
  signal blk00000003_sig000000d0 : STD_LOGIC; 
  signal blk00000003_sig000000cf : STD_LOGIC; 
  signal blk00000003_sig000000ce : STD_LOGIC; 
  signal blk00000003_sig000000cd : STD_LOGIC; 
  signal blk00000003_sig000000cc : STD_LOGIC; 
  signal blk00000003_sig000000cb : STD_LOGIC; 
  signal blk00000003_sig000000ca : STD_LOGIC; 
  signal blk00000003_sig000000c9 : STD_LOGIC; 
  signal blk00000003_sig000000c8 : STD_LOGIC; 
  signal blk00000003_sig000000c7 : STD_LOGIC; 
  signal blk00000003_sig000000c6 : STD_LOGIC; 
  signal blk00000003_sig000000c5 : STD_LOGIC; 
  signal blk00000003_sig000000c4 : STD_LOGIC; 
  signal blk00000003_sig000000c3 : STD_LOGIC; 
  signal blk00000003_sig000000c2 : STD_LOGIC; 
  signal blk00000003_sig000000c1 : STD_LOGIC; 
  signal blk00000003_sig000000c0 : STD_LOGIC; 
  signal blk00000003_sig000000bf : STD_LOGIC; 
  signal blk00000003_sig000000be : STD_LOGIC; 
  signal blk00000003_sig000000bd : STD_LOGIC; 
  signal blk00000003_sig000000bc : STD_LOGIC; 
  signal blk00000003_sig000000bb : STD_LOGIC; 
  signal blk00000003_sig000000ba : STD_LOGIC; 
  signal blk00000003_sig000000b9 : STD_LOGIC; 
  signal blk00000003_sig000000b8 : STD_LOGIC; 
  signal blk00000003_sig000000b7 : STD_LOGIC; 
  signal blk00000003_sig000000b6 : STD_LOGIC; 
  signal blk00000003_sig000000b5 : STD_LOGIC; 
  signal blk00000003_sig000000b4 : STD_LOGIC; 
  signal blk00000003_sig000000b3 : STD_LOGIC; 
  signal blk00000003_sig000000b2 : STD_LOGIC; 
  signal blk00000003_sig000000b1 : STD_LOGIC; 
  signal blk00000003_sig000000b0 : STD_LOGIC; 
  signal blk00000003_sig000000af : STD_LOGIC; 
  signal blk00000003_sig000000ae : STD_LOGIC; 
  signal blk00000003_sig000000ad : STD_LOGIC; 
  signal blk00000003_sig000000ac : STD_LOGIC; 
  signal blk00000003_sig000000ab : STD_LOGIC; 
  signal blk00000003_sig000000aa : STD_LOGIC; 
  signal blk00000003_sig000000a9 : STD_LOGIC; 
  signal blk00000003_sig000000a8 : STD_LOGIC; 
  signal blk00000003_sig000000a7 : STD_LOGIC; 
  signal blk00000003_sig000000a6 : STD_LOGIC; 
  signal blk00000003_sig000000a5 : STD_LOGIC; 
  signal blk00000003_sig000000a4 : STD_LOGIC; 
  signal blk00000003_sig000000a3 : STD_LOGIC; 
  signal blk00000003_sig000000a2 : STD_LOGIC; 
  signal blk00000003_sig000000a1 : STD_LOGIC; 
  signal blk00000003_sig000000a0 : STD_LOGIC; 
  signal blk00000003_sig0000009f : STD_LOGIC; 
  signal blk00000003_sig0000009e : STD_LOGIC; 
  signal blk00000003_sig0000009d : STD_LOGIC; 
  signal blk00000003_sig0000009c : STD_LOGIC; 
  signal blk00000003_sig0000009b : STD_LOGIC; 
  signal blk00000003_sig0000009a : STD_LOGIC; 
  signal blk00000003_sig00000099 : STD_LOGIC; 
  signal blk00000003_sig00000098 : STD_LOGIC; 
  signal blk00000003_sig00000097 : STD_LOGIC; 
  signal blk00000003_sig00000096 : STD_LOGIC; 
  signal blk00000003_sig00000095 : STD_LOGIC; 
  signal blk00000003_sig00000094 : STD_LOGIC; 
  signal blk00000003_sig00000093 : STD_LOGIC; 
  signal blk00000003_sig00000092 : STD_LOGIC; 
  signal blk00000003_sig00000091 : STD_LOGIC; 
  signal blk00000003_sig00000090 : STD_LOGIC; 
  signal blk00000003_sig0000008f : STD_LOGIC; 
  signal blk00000003_sig0000008e : STD_LOGIC; 
  signal blk00000003_sig0000008d : STD_LOGIC; 
  signal blk00000003_sig0000008c : STD_LOGIC; 
  signal blk00000003_sig0000008b : STD_LOGIC; 
  signal blk00000003_sig0000008a : STD_LOGIC; 
  signal blk00000003_sig00000089 : STD_LOGIC; 
  signal blk00000003_sig00000088 : STD_LOGIC; 
  signal blk00000003_sig00000087 : STD_LOGIC; 
  signal blk00000003_sig00000086 : STD_LOGIC; 
  signal blk00000003_sig00000085 : STD_LOGIC; 
  signal blk00000003_sig00000084 : STD_LOGIC; 
  signal blk00000003_sig00000083 : STD_LOGIC; 
  signal blk00000003_sig00000082 : STD_LOGIC; 
  signal blk00000003_sig00000081 : STD_LOGIC; 
  signal blk00000003_sig00000080 : STD_LOGIC; 
  signal blk00000003_sig0000007f : STD_LOGIC; 
  signal blk00000003_sig0000007e : STD_LOGIC; 
  signal blk00000003_sig0000007d : STD_LOGIC; 
  signal blk00000003_sig0000007c : STD_LOGIC; 
  signal blk00000003_sig0000007b : STD_LOGIC; 
  signal blk00000003_sig0000007a : STD_LOGIC; 
  signal blk00000003_sig00000079 : STD_LOGIC; 
  signal blk00000003_sig00000078 : STD_LOGIC; 
  signal blk00000003_sig00000077 : STD_LOGIC; 
  signal blk00000003_sig00000076 : STD_LOGIC; 
  signal blk00000003_sig00000075 : STD_LOGIC; 
  signal blk00000003_sig00000074 : STD_LOGIC; 
  signal blk00000003_sig00000073 : STD_LOGIC; 
  signal blk00000003_sig00000072 : STD_LOGIC; 
  signal blk00000003_sig00000071 : STD_LOGIC; 
  signal blk00000003_sig00000070 : STD_LOGIC; 
  signal blk00000003_sig0000006f : STD_LOGIC; 
  signal blk00000003_sig0000006e : STD_LOGIC; 
  signal blk00000003_sig0000006d : STD_LOGIC; 
  signal blk00000003_sig0000006c : STD_LOGIC; 
  signal blk00000003_sig0000006b : STD_LOGIC; 
  signal blk00000003_sig0000006a : STD_LOGIC; 
  signal blk00000003_sig00000069 : STD_LOGIC; 
  signal blk00000003_sig00000068 : STD_LOGIC; 
  signal blk00000003_sig00000067 : STD_LOGIC; 
  signal blk00000003_sig00000066 : STD_LOGIC; 
  signal blk00000003_sig00000065 : STD_LOGIC; 
  signal blk00000003_sig00000064 : STD_LOGIC; 
  signal blk00000003_sig00000063 : STD_LOGIC; 
  signal blk00000003_sig00000062 : STD_LOGIC; 
  signal blk00000003_sig00000061 : STD_LOGIC; 
  signal blk00000003_sig00000060 : STD_LOGIC; 
  signal blk00000003_sig0000005f : STD_LOGIC; 
  signal blk00000003_sig0000005e : STD_LOGIC; 
  signal blk00000003_sig0000005d : STD_LOGIC; 
  signal blk00000003_sig0000005c : STD_LOGIC; 
  signal blk00000003_sig0000005b : STD_LOGIC; 
  signal blk00000003_sig0000005a : STD_LOGIC; 
  signal blk00000003_sig00000059 : STD_LOGIC; 
  signal blk00000003_sig00000058 : STD_LOGIC; 
  signal blk00000003_sig00000057 : STD_LOGIC; 
  signal blk00000003_sig00000056 : STD_LOGIC; 
  signal blk00000003_sig00000055 : STD_LOGIC; 
  signal blk00000003_sig00000053 : STD_LOGIC; 
  signal NLW_blk00000001_P_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000002_G_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000003_blk00000186_O_UNCONNECTED : STD_LOGIC; 
begin
  rfd <= NlwRenamedSig_OI_rfd;
  blk00000001 : VCC
    port map (
      P => NLW_blk00000001_P_UNCONNECTED
    );
  blk00000002 : GND
    port map (
      G => NLW_blk00000002_G_UNCONNECTED
    );
  blk00000003_blk00000a38 : INV
    port map (
      I => blk00000003_sig000001db,
      O => blk00000003_sig000001e5
    );
  blk00000003_blk00000a37 : INV
    port map (
      I => blk00000003_sig000001dc,
      O => blk00000003_sig000001e8
    );
  blk00000003_blk00000a36 : INV
    port map (
      I => blk00000003_sig000001dd,
      O => blk00000003_sig000001eb
    );
  blk00000003_blk00000a35 : INV
    port map (
      I => blk00000003_sig000001de,
      O => blk00000003_sig000001ee
    );
  blk00000003_blk00000a34 : INV
    port map (
      I => blk00000003_sig000001df,
      O => blk00000003_sig000001f1
    );
  blk00000003_blk00000a33 : INV
    port map (
      I => blk00000003_sig000001e0,
      O => blk00000003_sig000001f4
    );
  blk00000003_blk00000a32 : INV
    port map (
      I => blk00000003_sig000001e1,
      O => blk00000003_sig000001f7
    );
  blk00000003_blk00000a31 : INV
    port map (
      I => blk00000003_sig00000a1b,
      O => blk00000003_sig0000009b
    );
  blk00000003_blk00000a30 : INV
    port map (
      I => blk00000003_sig00000a1c,
      O => blk00000003_sig0000009c
    );
  blk00000003_blk00000a2f : INV
    port map (
      I => blk00000003_sig00000a1d,
      O => blk00000003_sig0000009d
    );
  blk00000003_blk00000a2e : INV
    port map (
      I => blk00000003_sig00000a1e,
      O => blk00000003_sig0000009e
    );
  blk00000003_blk00000a2d : INV
    port map (
      I => blk00000003_sig00000a1f,
      O => blk00000003_sig0000009f
    );
  blk00000003_blk00000a2c : INV
    port map (
      I => blk00000003_sig00000a20,
      O => blk00000003_sig000000a0
    );
  blk00000003_blk00000a2b : INV
    port map (
      I => blk00000003_sig00000a21,
      O => blk00000003_sig000000a1
    );
  blk00000003_blk00000a2a : INV
    port map (
      I => blk00000003_sig00000a22,
      O => blk00000003_sig000000a2
    );
  blk00000003_blk00000a29 : INV
    port map (
      I => blk00000003_sig00000a23,
      O => blk00000003_sig000000a3
    );
  blk00000003_blk00000a28 : INV
    port map (
      I => blk00000003_sig00000a24,
      O => blk00000003_sig000000a4
    );
  blk00000003_blk00000a27 : INV
    port map (
      I => blk00000003_sig00000a25,
      O => blk00000003_sig000000a5
    );
  blk00000003_blk00000a26 : INV
    port map (
      I => blk00000003_sig00000a26,
      O => blk00000003_sig000000a6
    );
  blk00000003_blk00000a25 : INV
    port map (
      I => blk00000003_sig00000a27,
      O => blk00000003_sig000000a7
    );
  blk00000003_blk00000a24 : INV
    port map (
      I => blk00000003_sig00000a28,
      O => blk00000003_sig000000a8
    );
  blk00000003_blk00000a23 : INV
    port map (
      I => blk00000003_sig00000a29,
      O => blk00000003_sig000000a9
    );
  blk00000003_blk00000a22 : INV
    port map (
      I => blk00000003_sig00000a2a,
      O => blk00000003_sig000000aa
    );
  blk00000003_blk00000a21 : INV
    port map (
      I => blk00000003_sig00000a2b,
      O => blk00000003_sig000000ab
    );
  blk00000003_blk00000a20 : INV
    port map (
      I => blk00000003_sig00000a2c,
      O => blk00000003_sig000000ac
    );
  blk00000003_blk00000a1f : INV
    port map (
      I => blk00000003_sig00000a2d,
      O => blk00000003_sig000000ad
    );
  blk00000003_blk00000a1e : INV
    port map (
      I => blk00000003_sig00000a2e,
      O => blk00000003_sig000000ae
    );
  blk00000003_blk00000a1d : INV
    port map (
      I => blk00000003_sig00000a2f,
      O => blk00000003_sig000000af
    );
  blk00000003_blk00000a1c : INV
    port map (
      I => blk00000003_sig00000a30,
      O => blk00000003_sig000000b0
    );
  blk00000003_blk00000a1b : INV
    port map (
      I => blk00000003_sig00000a31,
      O => blk00000003_sig000000b1
    );
  blk00000003_blk00000a1a : INV
    port map (
      I => blk00000003_sig00000a32,
      O => blk00000003_sig000000b2
    );
  blk00000003_blk00000a19 : INV
    port map (
      I => blk00000003_sig00000a33,
      O => blk00000003_sig000000b3
    );
  blk00000003_blk00000a18 : INV
    port map (
      I => blk00000003_sig00000a34,
      O => blk00000003_sig000000b4
    );
  blk00000003_blk00000a17 : INV
    port map (
      I => blk00000003_sig00000a35,
      O => blk00000003_sig000000b5
    );
  blk00000003_blk00000a16 : INV
    port map (
      I => blk00000003_sig00000a36,
      O => blk00000003_sig000000b6
    );
  blk00000003_blk00000a15 : INV
    port map (
      I => blk00000003_sig00000a37,
      O => blk00000003_sig000000b7
    );
  blk00000003_blk00000a14 : INV
    port map (
      I => blk00000003_sig00000a38,
      O => blk00000003_sig000000b8
    );
  blk00000003_blk00000a13 : INV
    port map (
      I => blk00000003_sig00000a39,
      O => blk00000003_sig000000b9
    );
  blk00000003_blk00000a12 : INV
    port map (
      I => blk00000003_sig00000699,
      O => blk00000003_sig0000068c
    );
  blk00000003_blk00000a11 : INV
    port map (
      I => blk00000003_sig0000069a,
      O => blk00000003_sig00000667
    );
  blk00000003_blk00000a10 : INV
    port map (
      I => blk00000003_sig0000069b,
      O => blk00000003_sig00000642
    );
  blk00000003_blk00000a0f : INV
    port map (
      I => blk00000003_sig0000069c,
      O => blk00000003_sig0000061d
    );
  blk00000003_blk00000a0e : INV
    port map (
      I => blk00000003_sig0000069d,
      O => blk00000003_sig000005f8
    );
  blk00000003_blk00000a0d : INV
    port map (
      I => blk00000003_sig0000069e,
      O => blk00000003_sig000005d3
    );
  blk00000003_blk00000a0c : INV
    port map (
      I => blk00000003_sig0000069f,
      O => blk00000003_sig000005ae
    );
  blk00000003_blk00000a0b : INV
    port map (
      I => blk00000003_sig000006a0,
      O => blk00000003_sig00000588
    );
  blk00000003_blk00000a0a : INV
    port map (
      I => blk00000003_sig000006a1,
      O => blk00000003_sig00000562
    );
  blk00000003_blk00000a09 : INV
    port map (
      I => blk00000003_sig000006a2,
      O => blk00000003_sig0000053c
    );
  blk00000003_blk00000a08 : INV
    port map (
      I => blk00000003_sig000006a3,
      O => blk00000003_sig00000516
    );
  blk00000003_blk00000a07 : INV
    port map (
      I => blk00000003_sig000006a4,
      O => blk00000003_sig000004f0
    );
  blk00000003_blk00000a06 : INV
    port map (
      I => blk00000003_sig000006a5,
      O => blk00000003_sig000004ca
    );
  blk00000003_blk00000a05 : INV
    port map (
      I => blk00000003_sig000006a6,
      O => blk00000003_sig000004a4
    );
  blk00000003_blk00000a04 : INV
    port map (
      I => blk00000003_sig000006a7,
      O => blk00000003_sig0000047e
    );
  blk00000003_blk00000a03 : INV
    port map (
      I => blk00000003_sig000006a8,
      O => blk00000003_sig00000458
    );
  blk00000003_blk00000a02 : INV
    port map (
      I => blk00000003_sig000006a9,
      O => blk00000003_sig00000432
    );
  blk00000003_blk00000a01 : INV
    port map (
      I => blk00000003_sig000006aa,
      O => blk00000003_sig0000040c
    );
  blk00000003_blk00000a00 : INV
    port map (
      I => blk00000003_sig000006ab,
      O => blk00000003_sig000003e6
    );
  blk00000003_blk000009ff : INV
    port map (
      I => blk00000003_sig000006ac,
      O => blk00000003_sig000003c0
    );
  blk00000003_blk000009fe : INV
    port map (
      I => blk00000003_sig000006ad,
      O => blk00000003_sig0000039a
    );
  blk00000003_blk000009fd : INV
    port map (
      I => blk00000003_sig000006ae,
      O => blk00000003_sig00000374
    );
  blk00000003_blk000009fc : INV
    port map (
      I => blk00000003_sig000006af,
      O => blk00000003_sig0000034e
    );
  blk00000003_blk000009fb : INV
    port map (
      I => blk00000003_sig000006b0,
      O => blk00000003_sig00000328
    );
  blk00000003_blk000009fa : INV
    port map (
      I => blk00000003_sig00000077,
      O => blk00000003_sig00000302
    );
  blk00000003_blk000009f9 : INV
    port map (
      I => blk00000003_sig00000085,
      O => blk00000003_sig000002dc
    );
  blk00000003_blk000009f8 : INV
    port map (
      I => blk00000003_sig0000008b,
      O => blk00000003_sig000002b6
    );
  blk00000003_blk000009f7 : INV
    port map (
      I => blk00000003_sig00000090,
      O => blk00000003_sig00000290
    );
  blk00000003_blk000009f6 : INV
    port map (
      I => blk00000003_sig00000094,
      O => blk00000003_sig0000026a
    );
  blk00000003_blk000009f5 : INV
    port map (
      I => blk00000003_sig00000097,
      O => blk00000003_sig00000244
    );
  blk00000003_blk000009f4 : INV
    port map (
      I => blk00000003_sig00000099,
      O => blk00000003_sig0000021e
    );
  blk00000003_blk000009f3 : LUT1
    generic map(
      INIT => X"1"
    )
    port map (
      I0 => blk00000003_sig000001fc,
      O => blk00000003_sig00000099
    );
  blk00000003_blk000009f2 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000691,
      I1 => blk00000003_sig000000dc,
      I2 => blk00000003_sig00000690,
      O => blk00000003_sig00000a3b
    );
  blk00000003_blk000009f1 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000692,
      I1 => blk00000003_sig000000de,
      I2 => blk00000003_sig00000690,
      O => blk00000003_sig00000a3e
    );
  blk00000003_blk000009f0 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000693,
      I1 => blk00000003_sig000000e0,
      I2 => blk00000003_sig00000690,
      O => blk00000003_sig00000a41
    );
  blk00000003_blk000009ef : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000694,
      I1 => blk00000003_sig000000e2,
      I2 => blk00000003_sig00000690,
      O => blk00000003_sig00000a44
    );
  blk00000003_blk000009ee : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000695,
      I1 => blk00000003_sig000000e4,
      I2 => blk00000003_sig00000690,
      O => blk00000003_sig00000a47
    );
  blk00000003_blk000009ed : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000696,
      I1 => blk00000003_sig000000e6,
      I2 => blk00000003_sig00000690,
      O => blk00000003_sig00000a4a
    );
  blk00000003_blk000009ec : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000697,
      I1 => blk00000003_sig000000e8,
      I2 => blk00000003_sig00000690,
      O => blk00000003_sig00000a4d
    );
  blk00000003_blk000009eb : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000698,
      I1 => blk00000003_sig000000ea,
      I2 => blk00000003_sig00000690,
      O => blk00000003_sig00000a5a
    );
  blk00000003_blk000009ea : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000068a,
      I1 => blk00000003_sig00000699,
      O => blk00000003_sig0000066c
    );
  blk00000003_blk000009e9 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000683,
      I1 => blk00000003_sig000000db,
      I2 => blk00000003_sig00000699,
      O => blk00000003_sig0000066f
    );
  blk00000003_blk000009e8 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000684,
      I1 => blk00000003_sig000000dd,
      I2 => blk00000003_sig00000699,
      O => blk00000003_sig00000672
    );
  blk00000003_blk000009e7 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000685,
      I1 => blk00000003_sig000000df,
      I2 => blk00000003_sig00000699,
      O => blk00000003_sig00000675
    );
  blk00000003_blk000009e6 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000686,
      I1 => blk00000003_sig000000e1,
      I2 => blk00000003_sig00000699,
      O => blk00000003_sig00000678
    );
  blk00000003_blk000009e5 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000687,
      I1 => blk00000003_sig000000e3,
      I2 => blk00000003_sig00000699,
      O => blk00000003_sig0000067b
    );
  blk00000003_blk000009e4 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000688,
      I1 => blk00000003_sig000000e5,
      I2 => blk00000003_sig00000699,
      O => blk00000003_sig0000067e
    );
  blk00000003_blk000009e3 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000689,
      I1 => blk00000003_sig000000e7,
      I2 => blk00000003_sig00000699,
      O => blk00000003_sig00000681
    );
  blk00000003_blk000009e2 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000009a,
      I1 => blk00000003_sig000000e9,
      I2 => blk00000003_sig00000699,
      O => blk00000003_sig0000068d
    );
  blk00000003_blk000009e1 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000665,
      I1 => blk00000003_sig0000069a,
      O => blk00000003_sig00000647
    );
  blk00000003_blk000009e0 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000065e,
      I1 => blk00000003_sig000000eb,
      I2 => blk00000003_sig0000069a,
      O => blk00000003_sig0000064a
    );
  blk00000003_blk000009df : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000065f,
      I1 => blk00000003_sig000000ec,
      I2 => blk00000003_sig0000069a,
      O => blk00000003_sig0000064d
    );
  blk00000003_blk000009de : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000660,
      I1 => blk00000003_sig000000ed,
      I2 => blk00000003_sig0000069a,
      O => blk00000003_sig00000650
    );
  blk00000003_blk000009dd : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000661,
      I1 => blk00000003_sig000000ee,
      I2 => blk00000003_sig0000069a,
      O => blk00000003_sig00000653
    );
  blk00000003_blk000009dc : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000662,
      I1 => blk00000003_sig000000ef,
      I2 => blk00000003_sig0000069a,
      O => blk00000003_sig00000656
    );
  blk00000003_blk000009db : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000663,
      I1 => blk00000003_sig000000f0,
      I2 => blk00000003_sig0000069a,
      O => blk00000003_sig00000659
    );
  blk00000003_blk000009da : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000664,
      I1 => blk00000003_sig000000f1,
      I2 => blk00000003_sig0000069a,
      O => blk00000003_sig0000065c
    );
  blk00000003_blk000009d9 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000058,
      I1 => blk00000003_sig000000f2,
      I2 => blk00000003_sig0000069a,
      O => blk00000003_sig00000668
    );
  blk00000003_blk000009d8 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000640,
      I1 => blk00000003_sig0000069b,
      O => blk00000003_sig00000622
    );
  blk00000003_blk000009d7 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000639,
      I1 => blk00000003_sig000000f3,
      I2 => blk00000003_sig0000069b,
      O => blk00000003_sig00000625
    );
  blk00000003_blk000009d6 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000063a,
      I1 => blk00000003_sig000000f4,
      I2 => blk00000003_sig0000069b,
      O => blk00000003_sig00000628
    );
  blk00000003_blk000009d5 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000063b,
      I1 => blk00000003_sig000000f5,
      I2 => blk00000003_sig0000069b,
      O => blk00000003_sig0000062b
    );
  blk00000003_blk000009d4 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000063c,
      I1 => blk00000003_sig000000f6,
      I2 => blk00000003_sig0000069b,
      O => blk00000003_sig0000062e
    );
  blk00000003_blk000009d3 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000063d,
      I1 => blk00000003_sig000000f7,
      I2 => blk00000003_sig0000069b,
      O => blk00000003_sig00000631
    );
  blk00000003_blk000009d2 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000063e,
      I1 => blk00000003_sig000000f8,
      I2 => blk00000003_sig0000069b,
      O => blk00000003_sig00000634
    );
  blk00000003_blk000009d1 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000063f,
      I1 => blk00000003_sig000000f9,
      I2 => blk00000003_sig0000069b,
      O => blk00000003_sig00000637
    );
  blk00000003_blk000009d0 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000005c,
      I1 => blk00000003_sig000000fa,
      I2 => blk00000003_sig0000069b,
      O => blk00000003_sig00000643
    );
  blk00000003_blk000009cf : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000061b,
      I1 => blk00000003_sig0000069c,
      O => blk00000003_sig000005fd
    );
  blk00000003_blk000009ce : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000614,
      I1 => blk00000003_sig000000fb,
      I2 => blk00000003_sig0000069c,
      O => blk00000003_sig00000600
    );
  blk00000003_blk000009cd : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000615,
      I1 => blk00000003_sig000000fc,
      I2 => blk00000003_sig0000069c,
      O => blk00000003_sig00000603
    );
  blk00000003_blk000009cc : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000616,
      I1 => blk00000003_sig000000fd,
      I2 => blk00000003_sig0000069c,
      O => blk00000003_sig00000606
    );
  blk00000003_blk000009cb : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000617,
      I1 => blk00000003_sig000000fe,
      I2 => blk00000003_sig0000069c,
      O => blk00000003_sig00000609
    );
  blk00000003_blk000009ca : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000618,
      I1 => blk00000003_sig000000ff,
      I2 => blk00000003_sig0000069c,
      O => blk00000003_sig0000060c
    );
  blk00000003_blk000009c9 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000619,
      I1 => blk00000003_sig00000100,
      I2 => blk00000003_sig0000069c,
      O => blk00000003_sig0000060f
    );
  blk00000003_blk000009c8 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000061a,
      I1 => blk00000003_sig00000101,
      I2 => blk00000003_sig0000069c,
      O => blk00000003_sig00000612
    );
  blk00000003_blk000009c7 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000061,
      I1 => blk00000003_sig00000102,
      I2 => blk00000003_sig0000069c,
      O => blk00000003_sig0000061e
    );
  blk00000003_blk000009c6 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000005f6,
      I1 => blk00000003_sig0000069d,
      O => blk00000003_sig000005d8
    );
  blk00000003_blk000009c5 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005ef,
      I1 => blk00000003_sig00000103,
      I2 => blk00000003_sig0000069d,
      O => blk00000003_sig000005db
    );
  blk00000003_blk000009c4 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005f0,
      I1 => blk00000003_sig00000104,
      I2 => blk00000003_sig0000069d,
      O => blk00000003_sig000005de
    );
  blk00000003_blk000009c3 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005f1,
      I1 => blk00000003_sig00000105,
      I2 => blk00000003_sig0000069d,
      O => blk00000003_sig000005e1
    );
  blk00000003_blk000009c2 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005f2,
      I1 => blk00000003_sig00000106,
      I2 => blk00000003_sig0000069d,
      O => blk00000003_sig000005e4
    );
  blk00000003_blk000009c1 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005f3,
      I1 => blk00000003_sig00000107,
      I2 => blk00000003_sig0000069d,
      O => blk00000003_sig000005e7
    );
  blk00000003_blk000009c0 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005f4,
      I1 => blk00000003_sig00000108,
      I2 => blk00000003_sig0000069d,
      O => blk00000003_sig000005ea
    );
  blk00000003_blk000009bf : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005f5,
      I1 => blk00000003_sig00000109,
      I2 => blk00000003_sig0000069d,
      O => blk00000003_sig000005ed
    );
  blk00000003_blk000009be : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000067,
      I1 => blk00000003_sig0000010a,
      I2 => blk00000003_sig0000069d,
      O => blk00000003_sig000005f9
    );
  blk00000003_blk000009bd : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000005d1,
      I1 => blk00000003_sig0000069e,
      O => blk00000003_sig000005b3
    );
  blk00000003_blk000009bc : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005ca,
      I1 => blk00000003_sig0000010b,
      I2 => blk00000003_sig0000069e,
      O => blk00000003_sig000005b6
    );
  blk00000003_blk000009bb : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005cb,
      I1 => blk00000003_sig0000010c,
      I2 => blk00000003_sig0000069e,
      O => blk00000003_sig000005b9
    );
  blk00000003_blk000009ba : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005cc,
      I1 => blk00000003_sig0000010d,
      I2 => blk00000003_sig0000069e,
      O => blk00000003_sig000005bc
    );
  blk00000003_blk000009b9 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005cd,
      I1 => blk00000003_sig0000010e,
      I2 => blk00000003_sig0000069e,
      O => blk00000003_sig000005bf
    );
  blk00000003_blk000009b8 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005ce,
      I1 => blk00000003_sig0000010f,
      I2 => blk00000003_sig0000069e,
      O => blk00000003_sig000005c2
    );
  blk00000003_blk000009b7 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005cf,
      I1 => blk00000003_sig00000110,
      I2 => blk00000003_sig0000069e,
      O => blk00000003_sig000005c5
    );
  blk00000003_blk000009b6 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005d0,
      I1 => blk00000003_sig00000111,
      I2 => blk00000003_sig0000069e,
      O => blk00000003_sig000005c8
    );
  blk00000003_blk000009b5 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000006e,
      I1 => blk00000003_sig00000112,
      I2 => blk00000003_sig0000069e,
      O => blk00000003_sig000005d4
    );
  blk00000003_blk000009b4 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000005ac,
      I1 => blk00000003_sig0000069f,
      O => blk00000003_sig0000058e
    );
  blk00000003_blk000009b3 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005a5,
      I1 => blk00000003_sig00000113,
      I2 => blk00000003_sig0000069f,
      O => blk00000003_sig00000591
    );
  blk00000003_blk000009b2 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005a6,
      I1 => blk00000003_sig00000114,
      I2 => blk00000003_sig0000069f,
      O => blk00000003_sig00000594
    );
  blk00000003_blk000009b1 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005a7,
      I1 => blk00000003_sig00000115,
      I2 => blk00000003_sig0000069f,
      O => blk00000003_sig00000597
    );
  blk00000003_blk000009b0 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005a8,
      I1 => blk00000003_sig00000116,
      I2 => blk00000003_sig0000069f,
      O => blk00000003_sig0000059a
    );
  blk00000003_blk000009af : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005a9,
      I1 => blk00000003_sig00000117,
      I2 => blk00000003_sig0000069f,
      O => blk00000003_sig0000059d
    );
  blk00000003_blk000009ae : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005aa,
      I1 => blk00000003_sig00000118,
      I2 => blk00000003_sig0000069f,
      O => blk00000003_sig000005a0
    );
  blk00000003_blk000009ad : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000005ab,
      I1 => blk00000003_sig00000119,
      I2 => blk00000003_sig0000069f,
      O => blk00000003_sig000005a3
    );
  blk00000003_blk000009ac : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000076,
      I1 => blk00000003_sig0000011a,
      I2 => blk00000003_sig0000069f,
      O => blk00000003_sig000005af
    );
  blk00000003_blk000009ab : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000586,
      I1 => blk00000003_sig000006a0,
      O => blk00000003_sig00000568
    );
  blk00000003_blk000009aa : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000057f,
      I1 => blk00000003_sig0000011b,
      I2 => blk00000003_sig000006a0,
      O => blk00000003_sig0000056b
    );
  blk00000003_blk000009a9 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000580,
      I1 => blk00000003_sig0000011c,
      I2 => blk00000003_sig000006a0,
      O => blk00000003_sig0000056e
    );
  blk00000003_blk000009a8 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000581,
      I1 => blk00000003_sig0000011d,
      I2 => blk00000003_sig000006a0,
      O => blk00000003_sig00000571
    );
  blk00000003_blk000009a7 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000582,
      I1 => blk00000003_sig0000011e,
      I2 => blk00000003_sig000006a0,
      O => blk00000003_sig00000574
    );
  blk00000003_blk000009a6 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000583,
      I1 => blk00000003_sig0000011f,
      I2 => blk00000003_sig000006a0,
      O => blk00000003_sig00000577
    );
  blk00000003_blk000009a5 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000584,
      I1 => blk00000003_sig00000120,
      I2 => blk00000003_sig000006a0,
      O => blk00000003_sig0000057a
    );
  blk00000003_blk000009a4 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000585,
      I1 => blk00000003_sig00000121,
      I2 => blk00000003_sig000006a0,
      O => blk00000003_sig0000057d
    );
  blk00000003_blk000009a3 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000058b,
      I1 => blk00000003_sig00000122,
      I2 => blk00000003_sig000006a0,
      O => blk00000003_sig00000589
    );
  blk00000003_blk000009a2 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000560,
      I1 => blk00000003_sig000006a1,
      O => blk00000003_sig00000542
    );
  blk00000003_blk000009a1 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000559,
      I1 => blk00000003_sig00000123,
      I2 => blk00000003_sig000006a1,
      O => blk00000003_sig00000545
    );
  blk00000003_blk000009a0 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000055a,
      I1 => blk00000003_sig00000124,
      I2 => blk00000003_sig000006a1,
      O => blk00000003_sig00000548
    );
  blk00000003_blk0000099f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000055b,
      I1 => blk00000003_sig00000125,
      I2 => blk00000003_sig000006a1,
      O => blk00000003_sig0000054b
    );
  blk00000003_blk0000099e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000055c,
      I1 => blk00000003_sig00000126,
      I2 => blk00000003_sig000006a1,
      O => blk00000003_sig0000054e
    );
  blk00000003_blk0000099d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000055d,
      I1 => blk00000003_sig00000127,
      I2 => blk00000003_sig000006a1,
      O => blk00000003_sig00000551
    );
  blk00000003_blk0000099c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000055e,
      I1 => blk00000003_sig00000128,
      I2 => blk00000003_sig000006a1,
      O => blk00000003_sig00000554
    );
  blk00000003_blk0000099b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000055f,
      I1 => blk00000003_sig00000129,
      I2 => blk00000003_sig000006a1,
      O => blk00000003_sig00000557
    );
  blk00000003_blk0000099a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000565,
      I1 => blk00000003_sig0000012a,
      I2 => blk00000003_sig000006a1,
      O => blk00000003_sig00000563
    );
  blk00000003_blk00000999 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000053a,
      I1 => blk00000003_sig000006a2,
      O => blk00000003_sig0000051c
    );
  blk00000003_blk00000998 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000533,
      I1 => blk00000003_sig0000012b,
      I2 => blk00000003_sig000006a2,
      O => blk00000003_sig0000051f
    );
  blk00000003_blk00000997 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000534,
      I1 => blk00000003_sig0000012c,
      I2 => blk00000003_sig000006a2,
      O => blk00000003_sig00000522
    );
  blk00000003_blk00000996 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000535,
      I1 => blk00000003_sig0000012d,
      I2 => blk00000003_sig000006a2,
      O => blk00000003_sig00000525
    );
  blk00000003_blk00000995 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000536,
      I1 => blk00000003_sig0000012e,
      I2 => blk00000003_sig000006a2,
      O => blk00000003_sig00000528
    );
  blk00000003_blk00000994 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000537,
      I1 => blk00000003_sig0000012f,
      I2 => blk00000003_sig000006a2,
      O => blk00000003_sig0000052b
    );
  blk00000003_blk00000993 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000538,
      I1 => blk00000003_sig00000130,
      I2 => blk00000003_sig000006a2,
      O => blk00000003_sig0000052e
    );
  blk00000003_blk00000992 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000539,
      I1 => blk00000003_sig00000131,
      I2 => blk00000003_sig000006a2,
      O => blk00000003_sig00000531
    );
  blk00000003_blk00000991 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000053f,
      I1 => blk00000003_sig00000132,
      I2 => blk00000003_sig000006a2,
      O => blk00000003_sig0000053d
    );
  blk00000003_blk00000990 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000514,
      I1 => blk00000003_sig000006a3,
      O => blk00000003_sig000004f6
    );
  blk00000003_blk0000098f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000050d,
      I1 => blk00000003_sig00000133,
      I2 => blk00000003_sig000006a3,
      O => blk00000003_sig000004f9
    );
  blk00000003_blk0000098e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000050e,
      I1 => blk00000003_sig00000134,
      I2 => blk00000003_sig000006a3,
      O => blk00000003_sig000004fc
    );
  blk00000003_blk0000098d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000050f,
      I1 => blk00000003_sig00000135,
      I2 => blk00000003_sig000006a3,
      O => blk00000003_sig000004ff
    );
  blk00000003_blk0000098c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000510,
      I1 => blk00000003_sig00000136,
      I2 => blk00000003_sig000006a3,
      O => blk00000003_sig00000502
    );
  blk00000003_blk0000098b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000511,
      I1 => blk00000003_sig00000137,
      I2 => blk00000003_sig000006a3,
      O => blk00000003_sig00000505
    );
  blk00000003_blk0000098a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000512,
      I1 => blk00000003_sig00000138,
      I2 => blk00000003_sig000006a3,
      O => blk00000003_sig00000508
    );
  blk00000003_blk00000989 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000513,
      I1 => blk00000003_sig00000139,
      I2 => blk00000003_sig000006a3,
      O => blk00000003_sig0000050b
    );
  blk00000003_blk00000988 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000519,
      I1 => blk00000003_sig0000013a,
      I2 => blk00000003_sig000006a3,
      O => blk00000003_sig00000517
    );
  blk00000003_blk00000987 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000004ee,
      I1 => blk00000003_sig000006a4,
      O => blk00000003_sig000004d0
    );
  blk00000003_blk00000986 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004e7,
      I1 => blk00000003_sig0000013b,
      I2 => blk00000003_sig000006a4,
      O => blk00000003_sig000004d3
    );
  blk00000003_blk00000985 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004e8,
      I1 => blk00000003_sig0000013c,
      I2 => blk00000003_sig000006a4,
      O => blk00000003_sig000004d6
    );
  blk00000003_blk00000984 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004e9,
      I1 => blk00000003_sig0000013d,
      I2 => blk00000003_sig000006a4,
      O => blk00000003_sig000004d9
    );
  blk00000003_blk00000983 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004ea,
      I1 => blk00000003_sig0000013e,
      I2 => blk00000003_sig000006a4,
      O => blk00000003_sig000004dc
    );
  blk00000003_blk00000982 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004eb,
      I1 => blk00000003_sig0000013f,
      I2 => blk00000003_sig000006a4,
      O => blk00000003_sig000004df
    );
  blk00000003_blk00000981 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004ec,
      I1 => blk00000003_sig00000140,
      I2 => blk00000003_sig000006a4,
      O => blk00000003_sig000004e2
    );
  blk00000003_blk00000980 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004ed,
      I1 => blk00000003_sig00000141,
      I2 => blk00000003_sig000006a4,
      O => blk00000003_sig000004e5
    );
  blk00000003_blk0000097f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004f3,
      I1 => blk00000003_sig00000142,
      I2 => blk00000003_sig000006a4,
      O => blk00000003_sig000004f1
    );
  blk00000003_blk0000097e : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000004c8,
      I1 => blk00000003_sig000006a5,
      O => blk00000003_sig000004aa
    );
  blk00000003_blk0000097d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004c1,
      I1 => blk00000003_sig00000143,
      I2 => blk00000003_sig000006a5,
      O => blk00000003_sig000004ad
    );
  blk00000003_blk0000097c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004c2,
      I1 => blk00000003_sig00000144,
      I2 => blk00000003_sig000006a5,
      O => blk00000003_sig000004b0
    );
  blk00000003_blk0000097b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004c3,
      I1 => blk00000003_sig00000145,
      I2 => blk00000003_sig000006a5,
      O => blk00000003_sig000004b3
    );
  blk00000003_blk0000097a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004c4,
      I1 => blk00000003_sig00000146,
      I2 => blk00000003_sig000006a5,
      O => blk00000003_sig000004b6
    );
  blk00000003_blk00000979 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004c5,
      I1 => blk00000003_sig00000147,
      I2 => blk00000003_sig000006a5,
      O => blk00000003_sig000004b9
    );
  blk00000003_blk00000978 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004c6,
      I1 => blk00000003_sig00000148,
      I2 => blk00000003_sig000006a5,
      O => blk00000003_sig000004bc
    );
  blk00000003_blk00000977 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004c7,
      I1 => blk00000003_sig00000149,
      I2 => blk00000003_sig000006a5,
      O => blk00000003_sig000004bf
    );
  blk00000003_blk00000976 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004cd,
      I1 => blk00000003_sig0000014a,
      I2 => blk00000003_sig000006a5,
      O => blk00000003_sig000004cb
    );
  blk00000003_blk00000975 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000004a2,
      I1 => blk00000003_sig000006a6,
      O => blk00000003_sig00000484
    );
  blk00000003_blk00000974 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000049b,
      I1 => blk00000003_sig0000014b,
      I2 => blk00000003_sig000006a6,
      O => blk00000003_sig00000487
    );
  blk00000003_blk00000973 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000049c,
      I1 => blk00000003_sig0000014c,
      I2 => blk00000003_sig000006a6,
      O => blk00000003_sig0000048a
    );
  blk00000003_blk00000972 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000049d,
      I1 => blk00000003_sig0000014d,
      I2 => blk00000003_sig000006a6,
      O => blk00000003_sig0000048d
    );
  blk00000003_blk00000971 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000049e,
      I1 => blk00000003_sig0000014e,
      I2 => blk00000003_sig000006a6,
      O => blk00000003_sig00000490
    );
  blk00000003_blk00000970 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000049f,
      I1 => blk00000003_sig0000014f,
      I2 => blk00000003_sig000006a6,
      O => blk00000003_sig00000493
    );
  blk00000003_blk0000096f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004a0,
      I1 => blk00000003_sig00000150,
      I2 => blk00000003_sig000006a6,
      O => blk00000003_sig00000496
    );
  blk00000003_blk0000096e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004a1,
      I1 => blk00000003_sig00000151,
      I2 => blk00000003_sig000006a6,
      O => blk00000003_sig00000499
    );
  blk00000003_blk0000096d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004a7,
      I1 => blk00000003_sig00000152,
      I2 => blk00000003_sig000006a6,
      O => blk00000003_sig000004a5
    );
  blk00000003_blk0000096c : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000047c,
      I1 => blk00000003_sig000006a7,
      O => blk00000003_sig0000045e
    );
  blk00000003_blk0000096b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000475,
      I1 => blk00000003_sig00000153,
      I2 => blk00000003_sig000006a7,
      O => blk00000003_sig00000461
    );
  blk00000003_blk0000096a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000476,
      I1 => blk00000003_sig00000154,
      I2 => blk00000003_sig000006a7,
      O => blk00000003_sig00000464
    );
  blk00000003_blk00000969 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000477,
      I1 => blk00000003_sig00000155,
      I2 => blk00000003_sig000006a7,
      O => blk00000003_sig00000467
    );
  blk00000003_blk00000968 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000478,
      I1 => blk00000003_sig00000156,
      I2 => blk00000003_sig000006a7,
      O => blk00000003_sig0000046a
    );
  blk00000003_blk00000967 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000479,
      I1 => blk00000003_sig00000157,
      I2 => blk00000003_sig000006a7,
      O => blk00000003_sig0000046d
    );
  blk00000003_blk00000966 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000047a,
      I1 => blk00000003_sig00000158,
      I2 => blk00000003_sig000006a7,
      O => blk00000003_sig00000470
    );
  blk00000003_blk00000965 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000047b,
      I1 => blk00000003_sig00000159,
      I2 => blk00000003_sig000006a7,
      O => blk00000003_sig00000473
    );
  blk00000003_blk00000964 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000481,
      I1 => blk00000003_sig0000015a,
      I2 => blk00000003_sig000006a7,
      O => blk00000003_sig0000047f
    );
  blk00000003_blk00000963 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000456,
      I1 => blk00000003_sig000006a8,
      O => blk00000003_sig00000438
    );
  blk00000003_blk00000962 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000044f,
      I1 => blk00000003_sig0000015b,
      I2 => blk00000003_sig000006a8,
      O => blk00000003_sig0000043b
    );
  blk00000003_blk00000961 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000450,
      I1 => blk00000003_sig0000015c,
      I2 => blk00000003_sig000006a8,
      O => blk00000003_sig0000043e
    );
  blk00000003_blk00000960 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000451,
      I1 => blk00000003_sig0000015d,
      I2 => blk00000003_sig000006a8,
      O => blk00000003_sig00000441
    );
  blk00000003_blk0000095f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000452,
      I1 => blk00000003_sig0000015e,
      I2 => blk00000003_sig000006a8,
      O => blk00000003_sig00000444
    );
  blk00000003_blk0000095e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000453,
      I1 => blk00000003_sig0000015f,
      I2 => blk00000003_sig000006a8,
      O => blk00000003_sig00000447
    );
  blk00000003_blk0000095d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000454,
      I1 => blk00000003_sig00000160,
      I2 => blk00000003_sig000006a8,
      O => blk00000003_sig0000044a
    );
  blk00000003_blk0000095c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000455,
      I1 => blk00000003_sig00000161,
      I2 => blk00000003_sig000006a8,
      O => blk00000003_sig0000044d
    );
  blk00000003_blk0000095b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000045b,
      I1 => blk00000003_sig00000162,
      I2 => blk00000003_sig000006a8,
      O => blk00000003_sig00000459
    );
  blk00000003_blk0000095a : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000430,
      I1 => blk00000003_sig000006a9,
      O => blk00000003_sig00000412
    );
  blk00000003_blk00000959 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000429,
      I1 => blk00000003_sig00000163,
      I2 => blk00000003_sig000006a9,
      O => blk00000003_sig00000415
    );
  blk00000003_blk00000958 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000042a,
      I1 => blk00000003_sig00000164,
      I2 => blk00000003_sig000006a9,
      O => blk00000003_sig00000418
    );
  blk00000003_blk00000957 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000042b,
      I1 => blk00000003_sig00000165,
      I2 => blk00000003_sig000006a9,
      O => blk00000003_sig0000041b
    );
  blk00000003_blk00000956 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000042c,
      I1 => blk00000003_sig00000166,
      I2 => blk00000003_sig000006a9,
      O => blk00000003_sig0000041e
    );
  blk00000003_blk00000955 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000042d,
      I1 => blk00000003_sig00000167,
      I2 => blk00000003_sig000006a9,
      O => blk00000003_sig00000421
    );
  blk00000003_blk00000954 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000042e,
      I1 => blk00000003_sig00000168,
      I2 => blk00000003_sig000006a9,
      O => blk00000003_sig00000424
    );
  blk00000003_blk00000953 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000042f,
      I1 => blk00000003_sig00000169,
      I2 => blk00000003_sig000006a9,
      O => blk00000003_sig00000427
    );
  blk00000003_blk00000952 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000435,
      I1 => blk00000003_sig0000016a,
      I2 => blk00000003_sig000006a9,
      O => blk00000003_sig00000433
    );
  blk00000003_blk00000951 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000040a,
      I1 => blk00000003_sig000006aa,
      O => blk00000003_sig000003ec
    );
  blk00000003_blk00000950 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000403,
      I1 => blk00000003_sig0000016b,
      I2 => blk00000003_sig000006aa,
      O => blk00000003_sig000003ef
    );
  blk00000003_blk0000094f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000404,
      I1 => blk00000003_sig0000016c,
      I2 => blk00000003_sig000006aa,
      O => blk00000003_sig000003f2
    );
  blk00000003_blk0000094e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000405,
      I1 => blk00000003_sig0000016d,
      I2 => blk00000003_sig000006aa,
      O => blk00000003_sig000003f5
    );
  blk00000003_blk0000094d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000406,
      I1 => blk00000003_sig0000016e,
      I2 => blk00000003_sig000006aa,
      O => blk00000003_sig000003f8
    );
  blk00000003_blk0000094c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000407,
      I1 => blk00000003_sig0000016f,
      I2 => blk00000003_sig000006aa,
      O => blk00000003_sig000003fb
    );
  blk00000003_blk0000094b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000408,
      I1 => blk00000003_sig00000170,
      I2 => blk00000003_sig000006aa,
      O => blk00000003_sig000003fe
    );
  blk00000003_blk0000094a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000409,
      I1 => blk00000003_sig00000171,
      I2 => blk00000003_sig000006aa,
      O => blk00000003_sig00000401
    );
  blk00000003_blk00000949 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000040f,
      I1 => blk00000003_sig00000172,
      I2 => blk00000003_sig000006aa,
      O => blk00000003_sig0000040d
    );
  blk00000003_blk00000948 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000003e4,
      I1 => blk00000003_sig000006ab,
      O => blk00000003_sig000003c6
    );
  blk00000003_blk00000947 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003dd,
      I1 => blk00000003_sig00000173,
      I2 => blk00000003_sig000006ab,
      O => blk00000003_sig000003c9
    );
  blk00000003_blk00000946 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003de,
      I1 => blk00000003_sig00000174,
      I2 => blk00000003_sig000006ab,
      O => blk00000003_sig000003cc
    );
  blk00000003_blk00000945 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003df,
      I1 => blk00000003_sig00000175,
      I2 => blk00000003_sig000006ab,
      O => blk00000003_sig000003cf
    );
  blk00000003_blk00000944 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003e0,
      I1 => blk00000003_sig00000176,
      I2 => blk00000003_sig000006ab,
      O => blk00000003_sig000003d2
    );
  blk00000003_blk00000943 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003e1,
      I1 => blk00000003_sig00000177,
      I2 => blk00000003_sig000006ab,
      O => blk00000003_sig000003d5
    );
  blk00000003_blk00000942 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003e2,
      I1 => blk00000003_sig00000178,
      I2 => blk00000003_sig000006ab,
      O => blk00000003_sig000003d8
    );
  blk00000003_blk00000941 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003e3,
      I1 => blk00000003_sig00000179,
      I2 => blk00000003_sig000006ab,
      O => blk00000003_sig000003db
    );
  blk00000003_blk00000940 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003e9,
      I1 => blk00000003_sig0000017a,
      I2 => blk00000003_sig000006ab,
      O => blk00000003_sig000003e7
    );
  blk00000003_blk0000093f : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000003be,
      I1 => blk00000003_sig000006ac,
      O => blk00000003_sig000003a0
    );
  blk00000003_blk0000093e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003b7,
      I1 => blk00000003_sig0000017b,
      I2 => blk00000003_sig000006ac,
      O => blk00000003_sig000003a3
    );
  blk00000003_blk0000093d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003b8,
      I1 => blk00000003_sig0000017c,
      I2 => blk00000003_sig000006ac,
      O => blk00000003_sig000003a6
    );
  blk00000003_blk0000093c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003b9,
      I1 => blk00000003_sig0000017d,
      I2 => blk00000003_sig000006ac,
      O => blk00000003_sig000003a9
    );
  blk00000003_blk0000093b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003ba,
      I1 => blk00000003_sig0000017e,
      I2 => blk00000003_sig000006ac,
      O => blk00000003_sig000003ac
    );
  blk00000003_blk0000093a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003bb,
      I1 => blk00000003_sig0000017f,
      I2 => blk00000003_sig000006ac,
      O => blk00000003_sig000003af
    );
  blk00000003_blk00000939 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003bc,
      I1 => blk00000003_sig00000180,
      I2 => blk00000003_sig000006ac,
      O => blk00000003_sig000003b2
    );
  blk00000003_blk00000938 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003bd,
      I1 => blk00000003_sig00000181,
      I2 => blk00000003_sig000006ac,
      O => blk00000003_sig000003b5
    );
  blk00000003_blk00000937 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003c3,
      I1 => blk00000003_sig00000182,
      I2 => blk00000003_sig000006ac,
      O => blk00000003_sig000003c1
    );
  blk00000003_blk00000936 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000398,
      I1 => blk00000003_sig000006ad,
      O => blk00000003_sig0000037a
    );
  blk00000003_blk00000935 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000391,
      I1 => blk00000003_sig00000183,
      I2 => blk00000003_sig000006ad,
      O => blk00000003_sig0000037d
    );
  blk00000003_blk00000934 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000392,
      I1 => blk00000003_sig00000184,
      I2 => blk00000003_sig000006ad,
      O => blk00000003_sig00000380
    );
  blk00000003_blk00000933 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000393,
      I1 => blk00000003_sig00000185,
      I2 => blk00000003_sig000006ad,
      O => blk00000003_sig00000383
    );
  blk00000003_blk00000932 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000394,
      I1 => blk00000003_sig00000186,
      I2 => blk00000003_sig000006ad,
      O => blk00000003_sig00000386
    );
  blk00000003_blk00000931 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000395,
      I1 => blk00000003_sig00000187,
      I2 => blk00000003_sig000006ad,
      O => blk00000003_sig00000389
    );
  blk00000003_blk00000930 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000396,
      I1 => blk00000003_sig00000188,
      I2 => blk00000003_sig000006ad,
      O => blk00000003_sig0000038c
    );
  blk00000003_blk0000092f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000397,
      I1 => blk00000003_sig00000189,
      I2 => blk00000003_sig000006ad,
      O => blk00000003_sig0000038f
    );
  blk00000003_blk0000092e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000039d,
      I1 => blk00000003_sig0000018a,
      I2 => blk00000003_sig000006ad,
      O => blk00000003_sig0000039b
    );
  blk00000003_blk0000092d : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000372,
      I1 => blk00000003_sig000006ae,
      O => blk00000003_sig00000354
    );
  blk00000003_blk0000092c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000036b,
      I1 => blk00000003_sig0000018b,
      I2 => blk00000003_sig000006ae,
      O => blk00000003_sig00000357
    );
  blk00000003_blk0000092b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000036c,
      I1 => blk00000003_sig0000018c,
      I2 => blk00000003_sig000006ae,
      O => blk00000003_sig0000035a
    );
  blk00000003_blk0000092a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000036d,
      I1 => blk00000003_sig0000018d,
      I2 => blk00000003_sig000006ae,
      O => blk00000003_sig0000035d
    );
  blk00000003_blk00000929 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000036e,
      I1 => blk00000003_sig0000018e,
      I2 => blk00000003_sig000006ae,
      O => blk00000003_sig00000360
    );
  blk00000003_blk00000928 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000036f,
      I1 => blk00000003_sig0000018f,
      I2 => blk00000003_sig000006ae,
      O => blk00000003_sig00000363
    );
  blk00000003_blk00000927 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000370,
      I1 => blk00000003_sig00000190,
      I2 => blk00000003_sig000006ae,
      O => blk00000003_sig00000366
    );
  blk00000003_blk00000926 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000371,
      I1 => blk00000003_sig00000191,
      I2 => blk00000003_sig000006ae,
      O => blk00000003_sig00000369
    );
  blk00000003_blk00000925 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000377,
      I1 => blk00000003_sig00000192,
      I2 => blk00000003_sig000006ae,
      O => blk00000003_sig00000375
    );
  blk00000003_blk00000924 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000034c,
      I1 => blk00000003_sig000006af,
      O => blk00000003_sig0000032e
    );
  blk00000003_blk00000923 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000345,
      I1 => blk00000003_sig00000193,
      I2 => blk00000003_sig000006af,
      O => blk00000003_sig00000331
    );
  blk00000003_blk00000922 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000346,
      I1 => blk00000003_sig00000194,
      I2 => blk00000003_sig000006af,
      O => blk00000003_sig00000334
    );
  blk00000003_blk00000921 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000347,
      I1 => blk00000003_sig00000195,
      I2 => blk00000003_sig000006af,
      O => blk00000003_sig00000337
    );
  blk00000003_blk00000920 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000348,
      I1 => blk00000003_sig00000196,
      I2 => blk00000003_sig000006af,
      O => blk00000003_sig0000033a
    );
  blk00000003_blk0000091f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000349,
      I1 => blk00000003_sig00000197,
      I2 => blk00000003_sig000006af,
      O => blk00000003_sig0000033d
    );
  blk00000003_blk0000091e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000034a,
      I1 => blk00000003_sig00000198,
      I2 => blk00000003_sig000006af,
      O => blk00000003_sig00000340
    );
  blk00000003_blk0000091d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000034b,
      I1 => blk00000003_sig00000199,
      I2 => blk00000003_sig000006af,
      O => blk00000003_sig00000343
    );
  blk00000003_blk0000091c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000351,
      I1 => blk00000003_sig0000019a,
      I2 => blk00000003_sig000006af,
      O => blk00000003_sig0000034f
    );
  blk00000003_blk0000091b : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000326,
      I1 => blk00000003_sig000006b0,
      O => blk00000003_sig00000308
    );
  blk00000003_blk0000091a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000031f,
      I1 => blk00000003_sig0000019b,
      I2 => blk00000003_sig000006b0,
      O => blk00000003_sig0000030b
    );
  blk00000003_blk00000919 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000320,
      I1 => blk00000003_sig0000019c,
      I2 => blk00000003_sig000006b0,
      O => blk00000003_sig0000030e
    );
  blk00000003_blk00000918 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000321,
      I1 => blk00000003_sig0000019d,
      I2 => blk00000003_sig000006b0,
      O => blk00000003_sig00000311
    );
  blk00000003_blk00000917 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000322,
      I1 => blk00000003_sig0000019e,
      I2 => blk00000003_sig000006b0,
      O => blk00000003_sig00000314
    );
  blk00000003_blk00000916 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000323,
      I1 => blk00000003_sig0000019f,
      I2 => blk00000003_sig000006b0,
      O => blk00000003_sig00000317
    );
  blk00000003_blk00000915 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000324,
      I1 => blk00000003_sig000001a0,
      I2 => blk00000003_sig000006b0,
      O => blk00000003_sig0000031a
    );
  blk00000003_blk00000914 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000325,
      I1 => blk00000003_sig000001a1,
      I2 => blk00000003_sig000006b0,
      O => blk00000003_sig0000031d
    );
  blk00000003_blk00000913 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000032b,
      I1 => blk00000003_sig000001a2,
      I2 => blk00000003_sig000006b0,
      O => blk00000003_sig00000329
    );
  blk00000003_blk00000912 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000300,
      I1 => blk00000003_sig00000077,
      O => blk00000003_sig000002e2
    );
  blk00000003_blk00000911 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002f9,
      I1 => blk00000003_sig000001a3,
      I2 => blk00000003_sig00000077,
      O => blk00000003_sig000002e5
    );
  blk00000003_blk00000910 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002fa,
      I1 => blk00000003_sig000001a4,
      I2 => blk00000003_sig00000077,
      O => blk00000003_sig000002e8
    );
  blk00000003_blk0000090f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002fb,
      I1 => blk00000003_sig000001a5,
      I2 => blk00000003_sig00000077,
      O => blk00000003_sig000002eb
    );
  blk00000003_blk0000090e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002fc,
      I1 => blk00000003_sig000001a6,
      I2 => blk00000003_sig00000077,
      O => blk00000003_sig000002ee
    );
  blk00000003_blk0000090d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002fd,
      I1 => blk00000003_sig000001a7,
      I2 => blk00000003_sig00000077,
      O => blk00000003_sig000002f1
    );
  blk00000003_blk0000090c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002fe,
      I1 => blk00000003_sig000001a8,
      I2 => blk00000003_sig00000077,
      O => blk00000003_sig000002f4
    );
  blk00000003_blk0000090b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002ff,
      I1 => blk00000003_sig000001a9,
      I2 => blk00000003_sig00000077,
      O => blk00000003_sig000002f7
    );
  blk00000003_blk0000090a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000305,
      I1 => blk00000003_sig000001aa,
      I2 => blk00000003_sig00000077,
      O => blk00000003_sig00000303
    );
  blk00000003_blk00000909 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000002da,
      I1 => blk00000003_sig00000085,
      O => blk00000003_sig000002bc
    );
  blk00000003_blk00000908 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002d3,
      I1 => blk00000003_sig000001ab,
      I2 => blk00000003_sig00000085,
      O => blk00000003_sig000002bf
    );
  blk00000003_blk00000907 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002d4,
      I1 => blk00000003_sig000001ac,
      I2 => blk00000003_sig00000085,
      O => blk00000003_sig000002c2
    );
  blk00000003_blk00000906 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002d5,
      I1 => blk00000003_sig000001ad,
      I2 => blk00000003_sig00000085,
      O => blk00000003_sig000002c5
    );
  blk00000003_blk00000905 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002d6,
      I1 => blk00000003_sig000001ae,
      I2 => blk00000003_sig00000085,
      O => blk00000003_sig000002c8
    );
  blk00000003_blk00000904 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002d7,
      I1 => blk00000003_sig000001af,
      I2 => blk00000003_sig00000085,
      O => blk00000003_sig000002cb
    );
  blk00000003_blk00000903 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002d8,
      I1 => blk00000003_sig000001b0,
      I2 => blk00000003_sig00000085,
      O => blk00000003_sig000002ce
    );
  blk00000003_blk00000902 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002d9,
      I1 => blk00000003_sig000001b1,
      I2 => blk00000003_sig00000085,
      O => blk00000003_sig000002d1
    );
  blk00000003_blk00000901 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002df,
      I1 => blk00000003_sig000001b2,
      I2 => blk00000003_sig00000085,
      O => blk00000003_sig000002dd
    );
  blk00000003_blk00000900 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000002b4,
      I1 => blk00000003_sig0000008b,
      O => blk00000003_sig00000296
    );
  blk00000003_blk000008ff : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002ad,
      I1 => blk00000003_sig000001b3,
      I2 => blk00000003_sig0000008b,
      O => blk00000003_sig00000299
    );
  blk00000003_blk000008fe : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002ae,
      I1 => blk00000003_sig000001b4,
      I2 => blk00000003_sig0000008b,
      O => blk00000003_sig0000029c
    );
  blk00000003_blk000008fd : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002af,
      I1 => blk00000003_sig000001b5,
      I2 => blk00000003_sig0000008b,
      O => blk00000003_sig0000029f
    );
  blk00000003_blk000008fc : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002b0,
      I1 => blk00000003_sig000001b6,
      I2 => blk00000003_sig0000008b,
      O => blk00000003_sig000002a2
    );
  blk00000003_blk000008fb : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002b1,
      I1 => blk00000003_sig000001b7,
      I2 => blk00000003_sig0000008b,
      O => blk00000003_sig000002a5
    );
  blk00000003_blk000008fa : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002b2,
      I1 => blk00000003_sig000001b8,
      I2 => blk00000003_sig0000008b,
      O => blk00000003_sig000002a8
    );
  blk00000003_blk000008f9 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002b3,
      I1 => blk00000003_sig000001b9,
      I2 => blk00000003_sig0000008b,
      O => blk00000003_sig000002ab
    );
  blk00000003_blk000008f8 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002b9,
      I1 => blk00000003_sig000001ba,
      I2 => blk00000003_sig0000008b,
      O => blk00000003_sig000002b7
    );
  blk00000003_blk000008f7 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000028e,
      I1 => blk00000003_sig00000090,
      O => blk00000003_sig00000270
    );
  blk00000003_blk000008f6 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000287,
      I1 => blk00000003_sig000001bb,
      I2 => blk00000003_sig00000090,
      O => blk00000003_sig00000273
    );
  blk00000003_blk000008f5 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000288,
      I1 => blk00000003_sig000001bc,
      I2 => blk00000003_sig00000090,
      O => blk00000003_sig00000276
    );
  blk00000003_blk000008f4 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000289,
      I1 => blk00000003_sig000001bd,
      I2 => blk00000003_sig00000090,
      O => blk00000003_sig00000279
    );
  blk00000003_blk000008f3 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000028a,
      I1 => blk00000003_sig000001be,
      I2 => blk00000003_sig00000090,
      O => blk00000003_sig0000027c
    );
  blk00000003_blk000008f2 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000028b,
      I1 => blk00000003_sig000001bf,
      I2 => blk00000003_sig00000090,
      O => blk00000003_sig0000027f
    );
  blk00000003_blk000008f1 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000028c,
      I1 => blk00000003_sig000001c0,
      I2 => blk00000003_sig00000090,
      O => blk00000003_sig00000282
    );
  blk00000003_blk000008f0 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000028d,
      I1 => blk00000003_sig000001c1,
      I2 => blk00000003_sig00000090,
      O => blk00000003_sig00000285
    );
  blk00000003_blk000008ef : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000293,
      I1 => blk00000003_sig000001c2,
      I2 => blk00000003_sig00000090,
      O => blk00000003_sig00000291
    );
  blk00000003_blk000008ee : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000268,
      I1 => blk00000003_sig00000094,
      O => blk00000003_sig0000024a
    );
  blk00000003_blk000008ed : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000261,
      I1 => blk00000003_sig000001c3,
      I2 => blk00000003_sig00000094,
      O => blk00000003_sig0000024d
    );
  blk00000003_blk000008ec : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000262,
      I1 => blk00000003_sig000001c4,
      I2 => blk00000003_sig00000094,
      O => blk00000003_sig00000250
    );
  blk00000003_blk000008eb : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000263,
      I1 => blk00000003_sig000001c5,
      I2 => blk00000003_sig00000094,
      O => blk00000003_sig00000253
    );
  blk00000003_blk000008ea : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000264,
      I1 => blk00000003_sig000001c6,
      I2 => blk00000003_sig00000094,
      O => blk00000003_sig00000256
    );
  blk00000003_blk000008e9 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000265,
      I1 => blk00000003_sig000001c7,
      I2 => blk00000003_sig00000094,
      O => blk00000003_sig00000259
    );
  blk00000003_blk000008e8 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000266,
      I1 => blk00000003_sig000001c8,
      I2 => blk00000003_sig00000094,
      O => blk00000003_sig0000025c
    );
  blk00000003_blk000008e7 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000267,
      I1 => blk00000003_sig000001c9,
      I2 => blk00000003_sig00000094,
      O => blk00000003_sig0000025f
    );
  blk00000003_blk000008e6 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000026d,
      I1 => blk00000003_sig000001ca,
      I2 => blk00000003_sig00000094,
      O => blk00000003_sig0000026b
    );
  blk00000003_blk000008e5 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000242,
      I1 => blk00000003_sig00000097,
      O => blk00000003_sig00000224
    );
  blk00000003_blk000008e4 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000023b,
      I1 => blk00000003_sig000001cb,
      I2 => blk00000003_sig00000097,
      O => blk00000003_sig00000227
    );
  blk00000003_blk000008e3 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000023c,
      I1 => blk00000003_sig000001cc,
      I2 => blk00000003_sig00000097,
      O => blk00000003_sig0000022a
    );
  blk00000003_blk000008e2 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000023d,
      I1 => blk00000003_sig000001cd,
      I2 => blk00000003_sig00000097,
      O => blk00000003_sig0000022d
    );
  blk00000003_blk000008e1 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000023e,
      I1 => blk00000003_sig000001ce,
      I2 => blk00000003_sig00000097,
      O => blk00000003_sig00000230
    );
  blk00000003_blk000008e0 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000023f,
      I1 => blk00000003_sig000001cf,
      I2 => blk00000003_sig00000097,
      O => blk00000003_sig00000233
    );
  blk00000003_blk000008df : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000240,
      I1 => blk00000003_sig000001d0,
      I2 => blk00000003_sig00000097,
      O => blk00000003_sig00000236
    );
  blk00000003_blk000008de : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000241,
      I1 => blk00000003_sig000001d1,
      I2 => blk00000003_sig00000097,
      O => blk00000003_sig00000239
    );
  blk00000003_blk000008dd : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000247,
      I1 => blk00000003_sig000001d2,
      I2 => blk00000003_sig00000097,
      O => blk00000003_sig00000245
    );
  blk00000003_blk000008dc : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000021c,
      I1 => blk00000003_sig00000099,
      O => blk00000003_sig000001fe
    );
  blk00000003_blk000008db : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000215,
      I1 => blk00000003_sig000001d3,
      I2 => blk00000003_sig00000099,
      O => blk00000003_sig00000201
    );
  blk00000003_blk000008da : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000216,
      I1 => blk00000003_sig000001d4,
      I2 => blk00000003_sig00000099,
      O => blk00000003_sig00000204
    );
  blk00000003_blk000008d9 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000217,
      I1 => blk00000003_sig000001d5,
      I2 => blk00000003_sig00000099,
      O => blk00000003_sig00000207
    );
  blk00000003_blk000008d8 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000218,
      I1 => blk00000003_sig000001d6,
      I2 => blk00000003_sig00000099,
      O => blk00000003_sig0000020a
    );
  blk00000003_blk000008d7 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000219,
      I1 => blk00000003_sig000001d7,
      I2 => blk00000003_sig00000099,
      O => blk00000003_sig0000020d
    );
  blk00000003_blk000008d6 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000021a,
      I1 => blk00000003_sig000001d8,
      I2 => blk00000003_sig00000099,
      O => blk00000003_sig00000210
    );
  blk00000003_blk000008d5 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000021b,
      I1 => blk00000003_sig000001d9,
      I2 => blk00000003_sig00000099,
      O => blk00000003_sig00000213
    );
  blk00000003_blk000008d4 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000221,
      I1 => blk00000003_sig000001da,
      I2 => blk00000003_sig00000099,
      O => blk00000003_sig0000021f
    );
  blk00000003_blk000008d3 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000000bb,
      I1 => blk00000003_sig000001e2,
      O => blk00000003_sig000001fa
    );
  blk00000003_blk000008d2 : LUT1
    generic map(
      INIT => X"1"
    )
    port map (
      I0 => blk00000003_sig00000690,
      O => blk00000003_sig000000ba
    );
  blk00000003_blk000008d1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a5b,
      Q => fractional(0)
    );
  blk00000003_blk000008d0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a4e,
      Q => fractional(1)
    );
  blk00000003_blk000008cf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a4b,
      Q => fractional(2)
    );
  blk00000003_blk000008ce : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a48,
      Q => fractional(3)
    );
  blk00000003_blk000008cd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a45,
      Q => fractional(4)
    );
  blk00000003_blk000008cc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a42,
      Q => fractional(5)
    );
  blk00000003_blk000008cb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a3f,
      Q => fractional(6)
    );
  blk00000003_blk000008ca : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a3c,
      Q => fractional(7)
    );
  blk00000003_blk000008c9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a50,
      Q => blk00000003_sig00000a5e
    );
  blk00000003_blk000008c8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a52,
      Q => blk00000003_sig00000a5d
    );
  blk00000003_blk000008c7 : MULT_AND
    port map (
      I0 => blk00000003_sig000000ea,
      I1 => blk00000003_sig00000690,
      LO => blk00000003_sig00000a5c
    );
  blk00000003_blk000008c6 : MULT_AND
    port map (
      I0 => blk00000003_sig000000e8,
      I1 => blk00000003_sig00000690,
      LO => blk00000003_sig00000a59
    );
  blk00000003_blk000008c5 : MULT_AND
    port map (
      I0 => blk00000003_sig000000e6,
      I1 => blk00000003_sig00000690,
      LO => blk00000003_sig00000a58
    );
  blk00000003_blk000008c4 : MULT_AND
    port map (
      I0 => blk00000003_sig000000e4,
      I1 => blk00000003_sig00000690,
      LO => blk00000003_sig00000a57
    );
  blk00000003_blk000008c3 : MULT_AND
    port map (
      I0 => blk00000003_sig000000e2,
      I1 => blk00000003_sig00000690,
      LO => blk00000003_sig00000a56
    );
  blk00000003_blk000008c2 : MULT_AND
    port map (
      I0 => blk00000003_sig000000e0,
      I1 => blk00000003_sig00000690,
      LO => blk00000003_sig00000a55
    );
  blk00000003_blk000008c1 : MULT_AND
    port map (
      I0 => blk00000003_sig000000de,
      I1 => blk00000003_sig00000690,
      LO => blk00000003_sig00000a54
    );
  blk00000003_blk000008c0 : MULT_AND
    port map (
      I0 => blk00000003_sig000000dc,
      I1 => blk00000003_sig00000690,
      LO => blk00000003_sig00000a53
    );
  blk00000003_blk000008bf : MULT_AND
    port map (
      I0 => blk00000003_sig00000053,
      I1 => blk00000003_sig00000690,
      LO => blk00000003_sig00000a51
    );
  blk00000003_blk000008be : MUXCY
    port map (
      CI => blk00000003_sig00000053,
      DI => blk00000003_sig00000a5c,
      S => blk00000003_sig00000a5a,
      O => blk00000003_sig00000a4c
    );
  blk00000003_blk000008bd : XORCY
    port map (
      CI => blk00000003_sig00000053,
      LI => blk00000003_sig00000a5a,
      O => blk00000003_sig00000a5b
    );
  blk00000003_blk000008bc : MUXCY
    port map (
      CI => blk00000003_sig00000a4c,
      DI => blk00000003_sig00000a59,
      S => blk00000003_sig00000a4d,
      O => blk00000003_sig00000a49
    );
  blk00000003_blk000008bb : MUXCY
    port map (
      CI => blk00000003_sig00000a49,
      DI => blk00000003_sig00000a58,
      S => blk00000003_sig00000a4a,
      O => blk00000003_sig00000a46
    );
  blk00000003_blk000008ba : MUXCY
    port map (
      CI => blk00000003_sig00000a46,
      DI => blk00000003_sig00000a57,
      S => blk00000003_sig00000a47,
      O => blk00000003_sig00000a43
    );
  blk00000003_blk000008b9 : MUXCY
    port map (
      CI => blk00000003_sig00000a43,
      DI => blk00000003_sig00000a56,
      S => blk00000003_sig00000a44,
      O => blk00000003_sig00000a40
    );
  blk00000003_blk000008b8 : MUXCY
    port map (
      CI => blk00000003_sig00000a40,
      DI => blk00000003_sig00000a55,
      S => blk00000003_sig00000a41,
      O => blk00000003_sig00000a3d
    );
  blk00000003_blk000008b7 : MUXCY
    port map (
      CI => blk00000003_sig00000a3d,
      DI => blk00000003_sig00000a54,
      S => blk00000003_sig00000a3e,
      O => blk00000003_sig00000a3a
    );
  blk00000003_blk000008b6 : MUXCY
    port map (
      CI => blk00000003_sig00000a3a,
      DI => blk00000003_sig00000a53,
      S => blk00000003_sig00000a3b,
      O => blk00000003_sig00000a4f
    );
  blk00000003_blk000008b5 : MUXCY
    port map (
      CI => blk00000003_sig00000a4f,
      DI => blk00000003_sig00000a51,
      S => blk00000003_sig00000053,
      O => blk00000003_sig00000a52
    );
  blk00000003_blk000008b4 : XORCY
    port map (
      CI => blk00000003_sig00000a4f,
      LI => blk00000003_sig00000053,
      O => blk00000003_sig00000a50
    );
  blk00000003_blk000008b3 : XORCY
    port map (
      CI => blk00000003_sig00000a4c,
      LI => blk00000003_sig00000a4d,
      O => blk00000003_sig00000a4e
    );
  blk00000003_blk000008b2 : XORCY
    port map (
      CI => blk00000003_sig00000a49,
      LI => blk00000003_sig00000a4a,
      O => blk00000003_sig00000a4b
    );
  blk00000003_blk000008b1 : XORCY
    port map (
      CI => blk00000003_sig00000a46,
      LI => blk00000003_sig00000a47,
      O => blk00000003_sig00000a48
    );
  blk00000003_blk000008b0 : XORCY
    port map (
      CI => blk00000003_sig00000a43,
      LI => blk00000003_sig00000a44,
      O => blk00000003_sig00000a45
    );
  blk00000003_blk000008af : XORCY
    port map (
      CI => blk00000003_sig00000a40,
      LI => blk00000003_sig00000a41,
      O => blk00000003_sig00000a42
    );
  blk00000003_blk000008ae : XORCY
    port map (
      CI => blk00000003_sig00000a3d,
      LI => blk00000003_sig00000a3e,
      O => blk00000003_sig00000a3f
    );
  blk00000003_blk000008ad : XORCY
    port map (
      CI => blk00000003_sig00000a3a,
      LI => blk00000003_sig00000a3b,
      O => blk00000003_sig00000a3c
    );
  blk00000003_blk000008ac : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000699,
      Q => blk00000003_sig00000a39
    );
  blk00000003_blk000008ab : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a1a,
      Q => blk00000003_sig00000a38
    );
  blk00000003_blk000008aa : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a19,
      Q => blk00000003_sig00000a37
    );
  blk00000003_blk000008a9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a18,
      Q => blk00000003_sig00000a36
    );
  blk00000003_blk000008a8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a17,
      Q => blk00000003_sig00000a35
    );
  blk00000003_blk000008a7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a16,
      Q => blk00000003_sig00000a34
    );
  blk00000003_blk000008a6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a15,
      Q => blk00000003_sig00000a33
    );
  blk00000003_blk000008a5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a14,
      Q => blk00000003_sig00000a32
    );
  blk00000003_blk000008a4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a13,
      Q => blk00000003_sig00000a31
    );
  blk00000003_blk000008a3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a12,
      Q => blk00000003_sig00000a30
    );
  blk00000003_blk000008a2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a11,
      Q => blk00000003_sig00000a2f
    );
  blk00000003_blk000008a1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a10,
      Q => blk00000003_sig00000a2e
    );
  blk00000003_blk000008a0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a0f,
      Q => blk00000003_sig00000a2d
    );
  blk00000003_blk0000089f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a0e,
      Q => blk00000003_sig00000a2c
    );
  blk00000003_blk0000089e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a0d,
      Q => blk00000003_sig00000a2b
    );
  blk00000003_blk0000089d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a0c,
      Q => blk00000003_sig00000a2a
    );
  blk00000003_blk0000089c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a0b,
      Q => blk00000003_sig00000a29
    );
  blk00000003_blk0000089b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a0a,
      Q => blk00000003_sig00000a28
    );
  blk00000003_blk0000089a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a09,
      Q => blk00000003_sig00000a27
    );
  blk00000003_blk00000899 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a08,
      Q => blk00000003_sig00000a26
    );
  blk00000003_blk00000898 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a07,
      Q => blk00000003_sig00000a25
    );
  blk00000003_blk00000897 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a06,
      Q => blk00000003_sig00000a24
    );
  blk00000003_blk00000896 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a05,
      Q => blk00000003_sig00000a23
    );
  blk00000003_blk00000895 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a04,
      Q => blk00000003_sig00000a22
    );
  blk00000003_blk00000894 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a03,
      Q => blk00000003_sig00000a21
    );
  blk00000003_blk00000893 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a02,
      Q => blk00000003_sig00000a20
    );
  blk00000003_blk00000892 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a01,
      Q => blk00000003_sig00000a1f
    );
  blk00000003_blk00000891 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000a00,
      Q => blk00000003_sig00000a1e
    );
  blk00000003_blk00000890 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009ff,
      Q => blk00000003_sig00000a1d
    );
  blk00000003_blk0000088f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009fe,
      Q => blk00000003_sig00000a1c
    );
  blk00000003_blk0000088e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009fd,
      Q => blk00000003_sig00000a1b
    );
  blk00000003_blk0000088d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000069a,
      Q => blk00000003_sig00000a1a
    );
  blk00000003_blk0000088c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009fc,
      Q => blk00000003_sig00000a19
    );
  blk00000003_blk0000088b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009fb,
      Q => blk00000003_sig00000a18
    );
  blk00000003_blk0000088a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009fa,
      Q => blk00000003_sig00000a17
    );
  blk00000003_blk00000889 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009f9,
      Q => blk00000003_sig00000a16
    );
  blk00000003_blk00000888 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009f8,
      Q => blk00000003_sig00000a15
    );
  blk00000003_blk00000887 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009f7,
      Q => blk00000003_sig00000a14
    );
  blk00000003_blk00000886 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009f6,
      Q => blk00000003_sig00000a13
    );
  blk00000003_blk00000885 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009f5,
      Q => blk00000003_sig00000a12
    );
  blk00000003_blk00000884 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009f4,
      Q => blk00000003_sig00000a11
    );
  blk00000003_blk00000883 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009f3,
      Q => blk00000003_sig00000a10
    );
  blk00000003_blk00000882 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009f2,
      Q => blk00000003_sig00000a0f
    );
  blk00000003_blk00000881 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009f1,
      Q => blk00000003_sig00000a0e
    );
  blk00000003_blk00000880 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009f0,
      Q => blk00000003_sig00000a0d
    );
  blk00000003_blk0000087f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009ef,
      Q => blk00000003_sig00000a0c
    );
  blk00000003_blk0000087e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009ee,
      Q => blk00000003_sig00000a0b
    );
  blk00000003_blk0000087d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009ed,
      Q => blk00000003_sig00000a0a
    );
  blk00000003_blk0000087c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009ec,
      Q => blk00000003_sig00000a09
    );
  blk00000003_blk0000087b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009eb,
      Q => blk00000003_sig00000a08
    );
  blk00000003_blk0000087a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009ea,
      Q => blk00000003_sig00000a07
    );
  blk00000003_blk00000879 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009e9,
      Q => blk00000003_sig00000a06
    );
  blk00000003_blk00000878 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009e8,
      Q => blk00000003_sig00000a05
    );
  blk00000003_blk00000877 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009e7,
      Q => blk00000003_sig00000a04
    );
  blk00000003_blk00000876 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009e6,
      Q => blk00000003_sig00000a03
    );
  blk00000003_blk00000875 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009e5,
      Q => blk00000003_sig00000a02
    );
  blk00000003_blk00000874 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009e4,
      Q => blk00000003_sig00000a01
    );
  blk00000003_blk00000873 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009e3,
      Q => blk00000003_sig00000a00
    );
  blk00000003_blk00000872 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009e2,
      Q => blk00000003_sig000009ff
    );
  blk00000003_blk00000871 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009e1,
      Q => blk00000003_sig000009fe
    );
  blk00000003_blk00000870 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009e0,
      Q => blk00000003_sig000009fd
    );
  blk00000003_blk0000086f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000069b,
      Q => blk00000003_sig000009fc
    );
  blk00000003_blk0000086e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009df,
      Q => blk00000003_sig000009fb
    );
  blk00000003_blk0000086d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009de,
      Q => blk00000003_sig000009fa
    );
  blk00000003_blk0000086c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009dd,
      Q => blk00000003_sig000009f9
    );
  blk00000003_blk0000086b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009dc,
      Q => blk00000003_sig000009f8
    );
  blk00000003_blk0000086a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009db,
      Q => blk00000003_sig000009f7
    );
  blk00000003_blk00000869 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009da,
      Q => blk00000003_sig000009f6
    );
  blk00000003_blk00000868 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009d9,
      Q => blk00000003_sig000009f5
    );
  blk00000003_blk00000867 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009d8,
      Q => blk00000003_sig000009f4
    );
  blk00000003_blk00000866 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009d7,
      Q => blk00000003_sig000009f3
    );
  blk00000003_blk00000865 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009d6,
      Q => blk00000003_sig000009f2
    );
  blk00000003_blk00000864 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009d5,
      Q => blk00000003_sig000009f1
    );
  blk00000003_blk00000863 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009d4,
      Q => blk00000003_sig000009f0
    );
  blk00000003_blk00000862 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009d3,
      Q => blk00000003_sig000009ef
    );
  blk00000003_blk00000861 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009d2,
      Q => blk00000003_sig000009ee
    );
  blk00000003_blk00000860 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009d1,
      Q => blk00000003_sig000009ed
    );
  blk00000003_blk0000085f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009d0,
      Q => blk00000003_sig000009ec
    );
  blk00000003_blk0000085e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009cf,
      Q => blk00000003_sig000009eb
    );
  blk00000003_blk0000085d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009ce,
      Q => blk00000003_sig000009ea
    );
  blk00000003_blk0000085c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009cd,
      Q => blk00000003_sig000009e9
    );
  blk00000003_blk0000085b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009cc,
      Q => blk00000003_sig000009e8
    );
  blk00000003_blk0000085a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009cb,
      Q => blk00000003_sig000009e7
    );
  blk00000003_blk00000859 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009ca,
      Q => blk00000003_sig000009e6
    );
  blk00000003_blk00000858 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009c9,
      Q => blk00000003_sig000009e5
    );
  blk00000003_blk00000857 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009c8,
      Q => blk00000003_sig000009e4
    );
  blk00000003_blk00000856 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009c7,
      Q => blk00000003_sig000009e3
    );
  blk00000003_blk00000855 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009c6,
      Q => blk00000003_sig000009e2
    );
  blk00000003_blk00000854 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009c5,
      Q => blk00000003_sig000009e1
    );
  blk00000003_blk00000853 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009c4,
      Q => blk00000003_sig000009e0
    );
  blk00000003_blk00000852 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000069c,
      Q => blk00000003_sig000009df
    );
  blk00000003_blk00000851 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009c3,
      Q => blk00000003_sig000009de
    );
  blk00000003_blk00000850 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009c2,
      Q => blk00000003_sig000009dd
    );
  blk00000003_blk0000084f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009c1,
      Q => blk00000003_sig000009dc
    );
  blk00000003_blk0000084e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009c0,
      Q => blk00000003_sig000009db
    );
  blk00000003_blk0000084d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009bf,
      Q => blk00000003_sig000009da
    );
  blk00000003_blk0000084c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009be,
      Q => blk00000003_sig000009d9
    );
  blk00000003_blk0000084b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009bd,
      Q => blk00000003_sig000009d8
    );
  blk00000003_blk0000084a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009bc,
      Q => blk00000003_sig000009d7
    );
  blk00000003_blk00000849 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009bb,
      Q => blk00000003_sig000009d6
    );
  blk00000003_blk00000848 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009ba,
      Q => blk00000003_sig000009d5
    );
  blk00000003_blk00000847 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009b9,
      Q => blk00000003_sig000009d4
    );
  blk00000003_blk00000846 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009b8,
      Q => blk00000003_sig000009d3
    );
  blk00000003_blk00000845 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009b7,
      Q => blk00000003_sig000009d2
    );
  blk00000003_blk00000844 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009b6,
      Q => blk00000003_sig000009d1
    );
  blk00000003_blk00000843 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009b5,
      Q => blk00000003_sig000009d0
    );
  blk00000003_blk00000842 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009b4,
      Q => blk00000003_sig000009cf
    );
  blk00000003_blk00000841 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009b3,
      Q => blk00000003_sig000009ce
    );
  blk00000003_blk00000840 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009b2,
      Q => blk00000003_sig000009cd
    );
  blk00000003_blk0000083f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009b1,
      Q => blk00000003_sig000009cc
    );
  blk00000003_blk0000083e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009b0,
      Q => blk00000003_sig000009cb
    );
  blk00000003_blk0000083d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009af,
      Q => blk00000003_sig000009ca
    );
  blk00000003_blk0000083c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009ae,
      Q => blk00000003_sig000009c9
    );
  blk00000003_blk0000083b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009ad,
      Q => blk00000003_sig000009c8
    );
  blk00000003_blk0000083a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009ac,
      Q => blk00000003_sig000009c7
    );
  blk00000003_blk00000839 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009ab,
      Q => blk00000003_sig000009c6
    );
  blk00000003_blk00000838 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009aa,
      Q => blk00000003_sig000009c5
    );
  blk00000003_blk00000837 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009a9,
      Q => blk00000003_sig000009c4
    );
  blk00000003_blk00000836 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000069d,
      Q => blk00000003_sig000009c3
    );
  blk00000003_blk00000835 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009a8,
      Q => blk00000003_sig000009c2
    );
  blk00000003_blk00000834 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009a7,
      Q => blk00000003_sig000009c1
    );
  blk00000003_blk00000833 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009a6,
      Q => blk00000003_sig000009c0
    );
  blk00000003_blk00000832 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009a5,
      Q => blk00000003_sig000009bf
    );
  blk00000003_blk00000831 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009a4,
      Q => blk00000003_sig000009be
    );
  blk00000003_blk00000830 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009a3,
      Q => blk00000003_sig000009bd
    );
  blk00000003_blk0000082f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009a2,
      Q => blk00000003_sig000009bc
    );
  blk00000003_blk0000082e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009a1,
      Q => blk00000003_sig000009bb
    );
  blk00000003_blk0000082d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000009a0,
      Q => blk00000003_sig000009ba
    );
  blk00000003_blk0000082c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000099f,
      Q => blk00000003_sig000009b9
    );
  blk00000003_blk0000082b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000099e,
      Q => blk00000003_sig000009b8
    );
  blk00000003_blk0000082a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000099d,
      Q => blk00000003_sig000009b7
    );
  blk00000003_blk00000829 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000099c,
      Q => blk00000003_sig000009b6
    );
  blk00000003_blk00000828 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000099b,
      Q => blk00000003_sig000009b5
    );
  blk00000003_blk00000827 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000099a,
      Q => blk00000003_sig000009b4
    );
  blk00000003_blk00000826 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000999,
      Q => blk00000003_sig000009b3
    );
  blk00000003_blk00000825 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000998,
      Q => blk00000003_sig000009b2
    );
  blk00000003_blk00000824 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000997,
      Q => blk00000003_sig000009b1
    );
  blk00000003_blk00000823 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000996,
      Q => blk00000003_sig000009b0
    );
  blk00000003_blk00000822 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000995,
      Q => blk00000003_sig000009af
    );
  blk00000003_blk00000821 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000994,
      Q => blk00000003_sig000009ae
    );
  blk00000003_blk00000820 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000993,
      Q => blk00000003_sig000009ad
    );
  blk00000003_blk0000081f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000992,
      Q => blk00000003_sig000009ac
    );
  blk00000003_blk0000081e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000991,
      Q => blk00000003_sig000009ab
    );
  blk00000003_blk0000081d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000990,
      Q => blk00000003_sig000009aa
    );
  blk00000003_blk0000081c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000098f,
      Q => blk00000003_sig000009a9
    );
  blk00000003_blk0000081b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000069e,
      Q => blk00000003_sig000009a8
    );
  blk00000003_blk0000081a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000098e,
      Q => blk00000003_sig000009a7
    );
  blk00000003_blk00000819 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000098d,
      Q => blk00000003_sig000009a6
    );
  blk00000003_blk00000818 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000098c,
      Q => blk00000003_sig000009a5
    );
  blk00000003_blk00000817 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000098b,
      Q => blk00000003_sig000009a4
    );
  blk00000003_blk00000816 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000098a,
      Q => blk00000003_sig000009a3
    );
  blk00000003_blk00000815 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000989,
      Q => blk00000003_sig000009a2
    );
  blk00000003_blk00000814 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000988,
      Q => blk00000003_sig000009a1
    );
  blk00000003_blk00000813 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000987,
      Q => blk00000003_sig000009a0
    );
  blk00000003_blk00000812 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000986,
      Q => blk00000003_sig0000099f
    );
  blk00000003_blk00000811 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000985,
      Q => blk00000003_sig0000099e
    );
  blk00000003_blk00000810 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000984,
      Q => blk00000003_sig0000099d
    );
  blk00000003_blk0000080f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000983,
      Q => blk00000003_sig0000099c
    );
  blk00000003_blk0000080e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000982,
      Q => blk00000003_sig0000099b
    );
  blk00000003_blk0000080d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000981,
      Q => blk00000003_sig0000099a
    );
  blk00000003_blk0000080c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000980,
      Q => blk00000003_sig00000999
    );
  blk00000003_blk0000080b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000097f,
      Q => blk00000003_sig00000998
    );
  blk00000003_blk0000080a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000097e,
      Q => blk00000003_sig00000997
    );
  blk00000003_blk00000809 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000097d,
      Q => blk00000003_sig00000996
    );
  blk00000003_blk00000808 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000097c,
      Q => blk00000003_sig00000995
    );
  blk00000003_blk00000807 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000097b,
      Q => blk00000003_sig00000994
    );
  blk00000003_blk00000806 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000097a,
      Q => blk00000003_sig00000993
    );
  blk00000003_blk00000805 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000979,
      Q => blk00000003_sig00000992
    );
  blk00000003_blk00000804 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000978,
      Q => blk00000003_sig00000991
    );
  blk00000003_blk00000803 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000977,
      Q => blk00000003_sig00000990
    );
  blk00000003_blk00000802 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000976,
      Q => blk00000003_sig0000098f
    );
  blk00000003_blk00000801 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000069f,
      Q => blk00000003_sig0000098e
    );
  blk00000003_blk00000800 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000975,
      Q => blk00000003_sig0000098d
    );
  blk00000003_blk000007ff : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000974,
      Q => blk00000003_sig0000098c
    );
  blk00000003_blk000007fe : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000973,
      Q => blk00000003_sig0000098b
    );
  blk00000003_blk000007fd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000972,
      Q => blk00000003_sig0000098a
    );
  blk00000003_blk000007fc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000971,
      Q => blk00000003_sig00000989
    );
  blk00000003_blk000007fb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000970,
      Q => blk00000003_sig00000988
    );
  blk00000003_blk000007fa : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000096f,
      Q => blk00000003_sig00000987
    );
  blk00000003_blk000007f9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000096e,
      Q => blk00000003_sig00000986
    );
  blk00000003_blk000007f8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000096d,
      Q => blk00000003_sig00000985
    );
  blk00000003_blk000007f7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000096c,
      Q => blk00000003_sig00000984
    );
  blk00000003_blk000007f6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000096b,
      Q => blk00000003_sig00000983
    );
  blk00000003_blk000007f5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000096a,
      Q => blk00000003_sig00000982
    );
  blk00000003_blk000007f4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000969,
      Q => blk00000003_sig00000981
    );
  blk00000003_blk000007f3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000968,
      Q => blk00000003_sig00000980
    );
  blk00000003_blk000007f2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000967,
      Q => blk00000003_sig0000097f
    );
  blk00000003_blk000007f1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000966,
      Q => blk00000003_sig0000097e
    );
  blk00000003_blk000007f0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000965,
      Q => blk00000003_sig0000097d
    );
  blk00000003_blk000007ef : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000964,
      Q => blk00000003_sig0000097c
    );
  blk00000003_blk000007ee : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000963,
      Q => blk00000003_sig0000097b
    );
  blk00000003_blk000007ed : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000962,
      Q => blk00000003_sig0000097a
    );
  blk00000003_blk000007ec : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000961,
      Q => blk00000003_sig00000979
    );
  blk00000003_blk000007eb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000960,
      Q => blk00000003_sig00000978
    );
  blk00000003_blk000007ea : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000095f,
      Q => blk00000003_sig00000977
    );
  blk00000003_blk000007e9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000095e,
      Q => blk00000003_sig00000976
    );
  blk00000003_blk000007e8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a0,
      Q => blk00000003_sig00000975
    );
  blk00000003_blk000007e7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000095d,
      Q => blk00000003_sig00000974
    );
  blk00000003_blk000007e6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000095c,
      Q => blk00000003_sig00000973
    );
  blk00000003_blk000007e5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000095b,
      Q => blk00000003_sig00000972
    );
  blk00000003_blk000007e4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000095a,
      Q => blk00000003_sig00000971
    );
  blk00000003_blk000007e3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000959,
      Q => blk00000003_sig00000970
    );
  blk00000003_blk000007e2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000958,
      Q => blk00000003_sig0000096f
    );
  blk00000003_blk000007e1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000957,
      Q => blk00000003_sig0000096e
    );
  blk00000003_blk000007e0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000956,
      Q => blk00000003_sig0000096d
    );
  blk00000003_blk000007df : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000955,
      Q => blk00000003_sig0000096c
    );
  blk00000003_blk000007de : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000954,
      Q => blk00000003_sig0000096b
    );
  blk00000003_blk000007dd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000953,
      Q => blk00000003_sig0000096a
    );
  blk00000003_blk000007dc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000952,
      Q => blk00000003_sig00000969
    );
  blk00000003_blk000007db : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000951,
      Q => blk00000003_sig00000968
    );
  blk00000003_blk000007da : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000950,
      Q => blk00000003_sig00000967
    );
  blk00000003_blk000007d9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000094f,
      Q => blk00000003_sig00000966
    );
  blk00000003_blk000007d8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000094e,
      Q => blk00000003_sig00000965
    );
  blk00000003_blk000007d7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000094d,
      Q => blk00000003_sig00000964
    );
  blk00000003_blk000007d6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000094c,
      Q => blk00000003_sig00000963
    );
  blk00000003_blk000007d5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000094b,
      Q => blk00000003_sig00000962
    );
  blk00000003_blk000007d4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000094a,
      Q => blk00000003_sig00000961
    );
  blk00000003_blk000007d3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000949,
      Q => blk00000003_sig00000960
    );
  blk00000003_blk000007d2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000948,
      Q => blk00000003_sig0000095f
    );
  blk00000003_blk000007d1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000947,
      Q => blk00000003_sig0000095e
    );
  blk00000003_blk000007d0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000946,
      Q => blk00000003_sig0000006f
    );
  blk00000003_blk000007cf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000945,
      Q => blk00000003_sig00000070
    );
  blk00000003_blk000007ce : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000944,
      Q => blk00000003_sig00000071
    );
  blk00000003_blk000007cd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000943,
      Q => blk00000003_sig00000072
    );
  blk00000003_blk000007cc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000942,
      Q => blk00000003_sig00000073
    );
  blk00000003_blk000007cb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000941,
      Q => blk00000003_sig00000074
    );
  blk00000003_blk000007ca : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000940,
      Q => blk00000003_sig00000075
    );
  blk00000003_blk000007c9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000093f,
      Q => blk00000003_sig0000058b
    );
  blk00000003_blk000007c8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a1,
      Q => blk00000003_sig0000095d
    );
  blk00000003_blk000007c7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000093e,
      Q => blk00000003_sig0000095c
    );
  blk00000003_blk000007c6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000093d,
      Q => blk00000003_sig0000095b
    );
  blk00000003_blk000007c5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000093c,
      Q => blk00000003_sig0000095a
    );
  blk00000003_blk000007c4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000093b,
      Q => blk00000003_sig00000959
    );
  blk00000003_blk000007c3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000093a,
      Q => blk00000003_sig00000958
    );
  blk00000003_blk000007c2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000939,
      Q => blk00000003_sig00000957
    );
  blk00000003_blk000007c1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000938,
      Q => blk00000003_sig00000956
    );
  blk00000003_blk000007c0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000937,
      Q => blk00000003_sig00000955
    );
  blk00000003_blk000007bf : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000936,
      Q => blk00000003_sig00000954
    );
  blk00000003_blk000007be : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000935,
      Q => blk00000003_sig00000953
    );
  blk00000003_blk000007bd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000934,
      Q => blk00000003_sig00000952
    );
  blk00000003_blk000007bc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000933,
      Q => blk00000003_sig00000951
    );
  blk00000003_blk000007bb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000932,
      Q => blk00000003_sig00000950
    );
  blk00000003_blk000007ba : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000931,
      Q => blk00000003_sig0000094f
    );
  blk00000003_blk000007b9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000930,
      Q => blk00000003_sig0000094e
    );
  blk00000003_blk000007b8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000092f,
      Q => blk00000003_sig0000094d
    );
  blk00000003_blk000007b7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000092e,
      Q => blk00000003_sig0000094c
    );
  blk00000003_blk000007b6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000092d,
      Q => blk00000003_sig0000094b
    );
  blk00000003_blk000007b5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000092c,
      Q => blk00000003_sig0000094a
    );
  blk00000003_blk000007b4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000092b,
      Q => blk00000003_sig00000949
    );
  blk00000003_blk000007b3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000092a,
      Q => blk00000003_sig00000948
    );
  blk00000003_blk000007b2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000929,
      Q => blk00000003_sig00000947
    );
  blk00000003_blk000007b1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000928,
      Q => blk00000003_sig00000946
    );
  blk00000003_blk000007b0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000927,
      Q => blk00000003_sig00000945
    );
  blk00000003_blk000007af : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000926,
      Q => blk00000003_sig00000944
    );
  blk00000003_blk000007ae : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000925,
      Q => blk00000003_sig00000943
    );
  blk00000003_blk000007ad : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000924,
      Q => blk00000003_sig00000942
    );
  blk00000003_blk000007ac : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000923,
      Q => blk00000003_sig00000941
    );
  blk00000003_blk000007ab : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000922,
      Q => blk00000003_sig00000940
    );
  blk00000003_blk000007aa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000921,
      Q => blk00000003_sig0000093f
    );
  blk00000003_blk000007a9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000920,
      Q => blk00000003_sig00000565
    );
  blk00000003_blk000007a8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a2,
      Q => blk00000003_sig0000093e
    );
  blk00000003_blk000007a7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000091f,
      Q => blk00000003_sig0000093d
    );
  blk00000003_blk000007a6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000091e,
      Q => blk00000003_sig0000093c
    );
  blk00000003_blk000007a5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000091d,
      Q => blk00000003_sig0000093b
    );
  blk00000003_blk000007a4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000091c,
      Q => blk00000003_sig0000093a
    );
  blk00000003_blk000007a3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000091b,
      Q => blk00000003_sig00000939
    );
  blk00000003_blk000007a2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000091a,
      Q => blk00000003_sig00000938
    );
  blk00000003_blk000007a1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000919,
      Q => blk00000003_sig00000937
    );
  blk00000003_blk000007a0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000918,
      Q => blk00000003_sig00000936
    );
  blk00000003_blk0000079f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000917,
      Q => blk00000003_sig00000935
    );
  blk00000003_blk0000079e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000916,
      Q => blk00000003_sig00000934
    );
  blk00000003_blk0000079d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000915,
      Q => blk00000003_sig00000933
    );
  blk00000003_blk0000079c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000914,
      Q => blk00000003_sig00000932
    );
  blk00000003_blk0000079b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000913,
      Q => blk00000003_sig00000931
    );
  blk00000003_blk0000079a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000912,
      Q => blk00000003_sig00000930
    );
  blk00000003_blk00000799 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000911,
      Q => blk00000003_sig0000092f
    );
  blk00000003_blk00000798 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000910,
      Q => blk00000003_sig0000092e
    );
  blk00000003_blk00000797 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000090f,
      Q => blk00000003_sig0000092d
    );
  blk00000003_blk00000796 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000090e,
      Q => blk00000003_sig0000092c
    );
  blk00000003_blk00000795 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000090d,
      Q => blk00000003_sig0000092b
    );
  blk00000003_blk00000794 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000090c,
      Q => blk00000003_sig0000092a
    );
  blk00000003_blk00000793 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000090b,
      Q => blk00000003_sig00000929
    );
  blk00000003_blk00000792 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000090a,
      Q => blk00000003_sig00000928
    );
  blk00000003_blk00000791 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000909,
      Q => blk00000003_sig00000927
    );
  blk00000003_blk00000790 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000908,
      Q => blk00000003_sig00000926
    );
  blk00000003_blk0000078f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000907,
      Q => blk00000003_sig00000925
    );
  blk00000003_blk0000078e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000906,
      Q => blk00000003_sig00000924
    );
  blk00000003_blk0000078d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000905,
      Q => blk00000003_sig00000923
    );
  blk00000003_blk0000078c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000904,
      Q => blk00000003_sig00000922
    );
  blk00000003_blk0000078b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000903,
      Q => blk00000003_sig00000921
    );
  blk00000003_blk0000078a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000902,
      Q => blk00000003_sig00000920
    );
  blk00000003_blk00000789 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000901,
      Q => blk00000003_sig0000053f
    );
  blk00000003_blk00000788 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a3,
      Q => blk00000003_sig0000091f
    );
  blk00000003_blk00000787 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000900,
      Q => blk00000003_sig0000091e
    );
  blk00000003_blk00000786 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008ff,
      Q => blk00000003_sig0000091d
    );
  blk00000003_blk00000785 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008fe,
      Q => blk00000003_sig0000091c
    );
  blk00000003_blk00000784 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008fd,
      Q => blk00000003_sig0000091b
    );
  blk00000003_blk00000783 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008fc,
      Q => blk00000003_sig0000091a
    );
  blk00000003_blk00000782 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008fb,
      Q => blk00000003_sig00000919
    );
  blk00000003_blk00000781 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008fa,
      Q => blk00000003_sig00000918
    );
  blk00000003_blk00000780 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008f9,
      Q => blk00000003_sig00000917
    );
  blk00000003_blk0000077f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008f8,
      Q => blk00000003_sig00000916
    );
  blk00000003_blk0000077e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008f7,
      Q => blk00000003_sig00000915
    );
  blk00000003_blk0000077d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008f6,
      Q => blk00000003_sig00000914
    );
  blk00000003_blk0000077c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008f5,
      Q => blk00000003_sig00000913
    );
  blk00000003_blk0000077b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008f4,
      Q => blk00000003_sig00000912
    );
  blk00000003_blk0000077a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008f3,
      Q => blk00000003_sig00000911
    );
  blk00000003_blk00000779 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008f2,
      Q => blk00000003_sig00000910
    );
  blk00000003_blk00000778 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008f1,
      Q => blk00000003_sig0000090f
    );
  blk00000003_blk00000777 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008f0,
      Q => blk00000003_sig0000090e
    );
  blk00000003_blk00000776 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008ef,
      Q => blk00000003_sig0000090d
    );
  blk00000003_blk00000775 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008ee,
      Q => blk00000003_sig0000090c
    );
  blk00000003_blk00000774 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008ed,
      Q => blk00000003_sig0000090b
    );
  blk00000003_blk00000773 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008ec,
      Q => blk00000003_sig0000090a
    );
  blk00000003_blk00000772 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008eb,
      Q => blk00000003_sig00000909
    );
  blk00000003_blk00000771 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008ea,
      Q => blk00000003_sig00000908
    );
  blk00000003_blk00000770 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008e9,
      Q => blk00000003_sig00000907
    );
  blk00000003_blk0000076f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008e8,
      Q => blk00000003_sig00000906
    );
  blk00000003_blk0000076e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008e7,
      Q => blk00000003_sig00000905
    );
  blk00000003_blk0000076d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008e6,
      Q => blk00000003_sig00000904
    );
  blk00000003_blk0000076c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008e5,
      Q => blk00000003_sig00000903
    );
  blk00000003_blk0000076b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008e4,
      Q => blk00000003_sig00000902
    );
  blk00000003_blk0000076a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008e3,
      Q => blk00000003_sig00000901
    );
  blk00000003_blk00000769 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008e2,
      Q => blk00000003_sig00000519
    );
  blk00000003_blk00000768 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a4,
      Q => blk00000003_sig00000900
    );
  blk00000003_blk00000767 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008e1,
      Q => blk00000003_sig000008ff
    );
  blk00000003_blk00000766 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008e0,
      Q => blk00000003_sig000008fe
    );
  blk00000003_blk00000765 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008df,
      Q => blk00000003_sig000008fd
    );
  blk00000003_blk00000764 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008de,
      Q => blk00000003_sig000008fc
    );
  blk00000003_blk00000763 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008dd,
      Q => blk00000003_sig000008fb
    );
  blk00000003_blk00000762 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008dc,
      Q => blk00000003_sig000008fa
    );
  blk00000003_blk00000761 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008db,
      Q => blk00000003_sig000008f9
    );
  blk00000003_blk00000760 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008da,
      Q => blk00000003_sig000008f8
    );
  blk00000003_blk0000075f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008d9,
      Q => blk00000003_sig000008f7
    );
  blk00000003_blk0000075e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008d8,
      Q => blk00000003_sig000008f6
    );
  blk00000003_blk0000075d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008d7,
      Q => blk00000003_sig000008f5
    );
  blk00000003_blk0000075c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008d6,
      Q => blk00000003_sig000008f4
    );
  blk00000003_blk0000075b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008d5,
      Q => blk00000003_sig000008f3
    );
  blk00000003_blk0000075a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008d4,
      Q => blk00000003_sig000008f2
    );
  blk00000003_blk00000759 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008d3,
      Q => blk00000003_sig000008f1
    );
  blk00000003_blk00000758 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008d2,
      Q => blk00000003_sig000008f0
    );
  blk00000003_blk00000757 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008d1,
      Q => blk00000003_sig000008ef
    );
  blk00000003_blk00000756 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008d0,
      Q => blk00000003_sig000008ee
    );
  blk00000003_blk00000755 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008cf,
      Q => blk00000003_sig000008ed
    );
  blk00000003_blk00000754 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008ce,
      Q => blk00000003_sig000008ec
    );
  blk00000003_blk00000753 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008cd,
      Q => blk00000003_sig000008eb
    );
  blk00000003_blk00000752 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008cc,
      Q => blk00000003_sig000008ea
    );
  blk00000003_blk00000751 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008cb,
      Q => blk00000003_sig000008e9
    );
  blk00000003_blk00000750 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008ca,
      Q => blk00000003_sig000008e8
    );
  blk00000003_blk0000074f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008c9,
      Q => blk00000003_sig000008e7
    );
  blk00000003_blk0000074e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008c8,
      Q => blk00000003_sig000008e6
    );
  blk00000003_blk0000074d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008c7,
      Q => blk00000003_sig000008e5
    );
  blk00000003_blk0000074c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008c6,
      Q => blk00000003_sig000008e4
    );
  blk00000003_blk0000074b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008c5,
      Q => blk00000003_sig000008e3
    );
  blk00000003_blk0000074a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008c4,
      Q => blk00000003_sig000008e2
    );
  blk00000003_blk00000749 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008c3,
      Q => blk00000003_sig000004f3
    );
  blk00000003_blk00000748 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a5,
      Q => blk00000003_sig000008e1
    );
  blk00000003_blk00000747 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008c2,
      Q => blk00000003_sig000008e0
    );
  blk00000003_blk00000746 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008c1,
      Q => blk00000003_sig000008df
    );
  blk00000003_blk00000745 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008c0,
      Q => blk00000003_sig000008de
    );
  blk00000003_blk00000744 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008bf,
      Q => blk00000003_sig000008dd
    );
  blk00000003_blk00000743 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008be,
      Q => blk00000003_sig000008dc
    );
  blk00000003_blk00000742 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008bd,
      Q => blk00000003_sig000008db
    );
  blk00000003_blk00000741 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008bc,
      Q => blk00000003_sig000008da
    );
  blk00000003_blk00000740 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008bb,
      Q => blk00000003_sig000008d9
    );
  blk00000003_blk0000073f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008ba,
      Q => blk00000003_sig000008d8
    );
  blk00000003_blk0000073e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008b9,
      Q => blk00000003_sig000008d7
    );
  blk00000003_blk0000073d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008b8,
      Q => blk00000003_sig000008d6
    );
  blk00000003_blk0000073c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008b7,
      Q => blk00000003_sig000008d5
    );
  blk00000003_blk0000073b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008b6,
      Q => blk00000003_sig000008d4
    );
  blk00000003_blk0000073a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008b5,
      Q => blk00000003_sig000008d3
    );
  blk00000003_blk00000739 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008b4,
      Q => blk00000003_sig000008d2
    );
  blk00000003_blk00000738 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008b3,
      Q => blk00000003_sig000008d1
    );
  blk00000003_blk00000737 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008b2,
      Q => blk00000003_sig000008d0
    );
  blk00000003_blk00000736 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008b1,
      Q => blk00000003_sig000008cf
    );
  blk00000003_blk00000735 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008b0,
      Q => blk00000003_sig000008ce
    );
  blk00000003_blk00000734 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008af,
      Q => blk00000003_sig000008cd
    );
  blk00000003_blk00000733 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008ae,
      Q => blk00000003_sig000008cc
    );
  blk00000003_blk00000732 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008ad,
      Q => blk00000003_sig000008cb
    );
  blk00000003_blk00000731 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008ac,
      Q => blk00000003_sig000008ca
    );
  blk00000003_blk00000730 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008ab,
      Q => blk00000003_sig000008c9
    );
  blk00000003_blk0000072f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008aa,
      Q => blk00000003_sig000008c8
    );
  blk00000003_blk0000072e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008a9,
      Q => blk00000003_sig000008c7
    );
  blk00000003_blk0000072d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008a8,
      Q => blk00000003_sig000008c6
    );
  blk00000003_blk0000072c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008a7,
      Q => blk00000003_sig000008c5
    );
  blk00000003_blk0000072b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008a6,
      Q => blk00000003_sig000008c4
    );
  blk00000003_blk0000072a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008a5,
      Q => blk00000003_sig000008c3
    );
  blk00000003_blk00000729 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008a4,
      Q => blk00000003_sig000004cd
    );
  blk00000003_blk00000728 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a6,
      Q => blk00000003_sig000008c2
    );
  blk00000003_blk00000727 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008a3,
      Q => blk00000003_sig000008c1
    );
  blk00000003_blk00000726 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008a2,
      Q => blk00000003_sig000008c0
    );
  blk00000003_blk00000725 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008a1,
      Q => blk00000003_sig000008bf
    );
  blk00000003_blk00000724 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008a0,
      Q => blk00000003_sig000008be
    );
  blk00000003_blk00000723 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000089f,
      Q => blk00000003_sig000008bd
    );
  blk00000003_blk00000722 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000089e,
      Q => blk00000003_sig000008bc
    );
  blk00000003_blk00000721 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000089d,
      Q => blk00000003_sig000008bb
    );
  blk00000003_blk00000720 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000089c,
      Q => blk00000003_sig000008ba
    );
  blk00000003_blk0000071f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000089b,
      Q => blk00000003_sig000008b9
    );
  blk00000003_blk0000071e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000089a,
      Q => blk00000003_sig000008b8
    );
  blk00000003_blk0000071d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000899,
      Q => blk00000003_sig000008b7
    );
  blk00000003_blk0000071c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000898,
      Q => blk00000003_sig000008b6
    );
  blk00000003_blk0000071b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000897,
      Q => blk00000003_sig000008b5
    );
  blk00000003_blk0000071a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000896,
      Q => blk00000003_sig000008b4
    );
  blk00000003_blk00000719 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000895,
      Q => blk00000003_sig000008b3
    );
  blk00000003_blk00000718 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000894,
      Q => blk00000003_sig000008b2
    );
  blk00000003_blk00000717 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000893,
      Q => blk00000003_sig000008b1
    );
  blk00000003_blk00000716 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000892,
      Q => blk00000003_sig000008b0
    );
  blk00000003_blk00000715 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000891,
      Q => blk00000003_sig000008af
    );
  blk00000003_blk00000714 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000890,
      Q => blk00000003_sig000008ae
    );
  blk00000003_blk00000713 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000088f,
      Q => blk00000003_sig000008ad
    );
  blk00000003_blk00000712 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000088e,
      Q => blk00000003_sig000008ac
    );
  blk00000003_blk00000711 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000088d,
      Q => blk00000003_sig000008ab
    );
  blk00000003_blk00000710 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000088c,
      Q => blk00000003_sig000008aa
    );
  blk00000003_blk0000070f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000088b,
      Q => blk00000003_sig000008a9
    );
  blk00000003_blk0000070e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000088a,
      Q => blk00000003_sig000008a8
    );
  blk00000003_blk0000070d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000889,
      Q => blk00000003_sig000008a7
    );
  blk00000003_blk0000070c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000888,
      Q => blk00000003_sig000008a6
    );
  blk00000003_blk0000070b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000887,
      Q => blk00000003_sig000008a5
    );
  blk00000003_blk0000070a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000886,
      Q => blk00000003_sig000008a4
    );
  blk00000003_blk00000709 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000885,
      Q => blk00000003_sig000004a7
    );
  blk00000003_blk00000708 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a7,
      Q => blk00000003_sig000008a3
    );
  blk00000003_blk00000707 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000884,
      Q => blk00000003_sig000008a2
    );
  blk00000003_blk00000706 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000883,
      Q => blk00000003_sig000008a1
    );
  blk00000003_blk00000705 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000882,
      Q => blk00000003_sig000008a0
    );
  blk00000003_blk00000704 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000881,
      Q => blk00000003_sig0000089f
    );
  blk00000003_blk00000703 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000880,
      Q => blk00000003_sig0000089e
    );
  blk00000003_blk00000702 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000087f,
      Q => blk00000003_sig0000089d
    );
  blk00000003_blk00000701 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000087e,
      Q => blk00000003_sig0000089c
    );
  blk00000003_blk00000700 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000087d,
      Q => blk00000003_sig0000089b
    );
  blk00000003_blk000006ff : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000087c,
      Q => blk00000003_sig0000089a
    );
  blk00000003_blk000006fe : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000087b,
      Q => blk00000003_sig00000899
    );
  blk00000003_blk000006fd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000087a,
      Q => blk00000003_sig00000898
    );
  blk00000003_blk000006fc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000879,
      Q => blk00000003_sig00000897
    );
  blk00000003_blk000006fb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000878,
      Q => blk00000003_sig00000896
    );
  blk00000003_blk000006fa : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000877,
      Q => blk00000003_sig00000895
    );
  blk00000003_blk000006f9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000876,
      Q => blk00000003_sig00000894
    );
  blk00000003_blk000006f8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000875,
      Q => blk00000003_sig00000893
    );
  blk00000003_blk000006f7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000874,
      Q => blk00000003_sig00000892
    );
  blk00000003_blk000006f6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000873,
      Q => blk00000003_sig00000891
    );
  blk00000003_blk000006f5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000872,
      Q => blk00000003_sig00000890
    );
  blk00000003_blk000006f4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000871,
      Q => blk00000003_sig0000088f
    );
  blk00000003_blk000006f3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000870,
      Q => blk00000003_sig0000088e
    );
  blk00000003_blk000006f2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000086f,
      Q => blk00000003_sig0000088d
    );
  blk00000003_blk000006f1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000086e,
      Q => blk00000003_sig0000088c
    );
  blk00000003_blk000006f0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000086d,
      Q => blk00000003_sig0000088b
    );
  blk00000003_blk000006ef : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000086c,
      Q => blk00000003_sig0000088a
    );
  blk00000003_blk000006ee : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000086b,
      Q => blk00000003_sig00000889
    );
  blk00000003_blk000006ed : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000086a,
      Q => blk00000003_sig00000888
    );
  blk00000003_blk000006ec : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000869,
      Q => blk00000003_sig00000887
    );
  blk00000003_blk000006eb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000868,
      Q => blk00000003_sig00000886
    );
  blk00000003_blk000006ea : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000867,
      Q => blk00000003_sig00000885
    );
  blk00000003_blk000006e9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000866,
      Q => blk00000003_sig00000481
    );
  blk00000003_blk000006e8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a8,
      Q => blk00000003_sig00000884
    );
  blk00000003_blk000006e7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000865,
      Q => blk00000003_sig00000883
    );
  blk00000003_blk000006e6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000864,
      Q => blk00000003_sig00000882
    );
  blk00000003_blk000006e5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000863,
      Q => blk00000003_sig00000881
    );
  blk00000003_blk000006e4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000862,
      Q => blk00000003_sig00000880
    );
  blk00000003_blk000006e3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000861,
      Q => blk00000003_sig0000087f
    );
  blk00000003_blk000006e2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000860,
      Q => blk00000003_sig0000087e
    );
  blk00000003_blk000006e1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000085f,
      Q => blk00000003_sig0000087d
    );
  blk00000003_blk000006e0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000085e,
      Q => blk00000003_sig0000087c
    );
  blk00000003_blk000006df : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000085d,
      Q => blk00000003_sig0000087b
    );
  blk00000003_blk000006de : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000085c,
      Q => blk00000003_sig0000087a
    );
  blk00000003_blk000006dd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000085b,
      Q => blk00000003_sig00000879
    );
  blk00000003_blk000006dc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000085a,
      Q => blk00000003_sig00000878
    );
  blk00000003_blk000006db : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000859,
      Q => blk00000003_sig00000877
    );
  blk00000003_blk000006da : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000858,
      Q => blk00000003_sig00000876
    );
  blk00000003_blk000006d9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000857,
      Q => blk00000003_sig00000875
    );
  blk00000003_blk000006d8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000856,
      Q => blk00000003_sig00000874
    );
  blk00000003_blk000006d7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000855,
      Q => blk00000003_sig00000873
    );
  blk00000003_blk000006d6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000854,
      Q => blk00000003_sig00000872
    );
  blk00000003_blk000006d5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000853,
      Q => blk00000003_sig00000871
    );
  blk00000003_blk000006d4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000852,
      Q => blk00000003_sig00000870
    );
  blk00000003_blk000006d3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000851,
      Q => blk00000003_sig0000086f
    );
  blk00000003_blk000006d2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000850,
      Q => blk00000003_sig0000086e
    );
  blk00000003_blk000006d1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000084f,
      Q => blk00000003_sig0000086d
    );
  blk00000003_blk000006d0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000084e,
      Q => blk00000003_sig0000086c
    );
  blk00000003_blk000006cf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000084d,
      Q => blk00000003_sig0000086b
    );
  blk00000003_blk000006ce : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000084c,
      Q => blk00000003_sig0000086a
    );
  blk00000003_blk000006cd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000084b,
      Q => blk00000003_sig00000869
    );
  blk00000003_blk000006cc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000084a,
      Q => blk00000003_sig00000868
    );
  blk00000003_blk000006cb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000849,
      Q => blk00000003_sig00000867
    );
  blk00000003_blk000006ca : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000848,
      Q => blk00000003_sig00000866
    );
  blk00000003_blk000006c9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000847,
      Q => blk00000003_sig0000045b
    );
  blk00000003_blk000006c8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a9,
      Q => blk00000003_sig00000865
    );
  blk00000003_blk000006c7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000846,
      Q => blk00000003_sig00000864
    );
  blk00000003_blk000006c6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000845,
      Q => blk00000003_sig00000863
    );
  blk00000003_blk000006c5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000844,
      Q => blk00000003_sig00000862
    );
  blk00000003_blk000006c4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000843,
      Q => blk00000003_sig00000861
    );
  blk00000003_blk000006c3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000842,
      Q => blk00000003_sig00000860
    );
  blk00000003_blk000006c2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000841,
      Q => blk00000003_sig0000085f
    );
  blk00000003_blk000006c1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000840,
      Q => blk00000003_sig0000085e
    );
  blk00000003_blk000006c0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000083f,
      Q => blk00000003_sig0000085d
    );
  blk00000003_blk000006bf : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000083e,
      Q => blk00000003_sig0000085c
    );
  blk00000003_blk000006be : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000083d,
      Q => blk00000003_sig0000085b
    );
  blk00000003_blk000006bd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000083c,
      Q => blk00000003_sig0000085a
    );
  blk00000003_blk000006bc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000083b,
      Q => blk00000003_sig00000859
    );
  blk00000003_blk000006bb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000083a,
      Q => blk00000003_sig00000858
    );
  blk00000003_blk000006ba : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000839,
      Q => blk00000003_sig00000857
    );
  blk00000003_blk000006b9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000838,
      Q => blk00000003_sig00000856
    );
  blk00000003_blk000006b8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000837,
      Q => blk00000003_sig00000855
    );
  blk00000003_blk000006b7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000836,
      Q => blk00000003_sig00000854
    );
  blk00000003_blk000006b6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000835,
      Q => blk00000003_sig00000853
    );
  blk00000003_blk000006b5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000834,
      Q => blk00000003_sig00000852
    );
  blk00000003_blk000006b4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000833,
      Q => blk00000003_sig00000851
    );
  blk00000003_blk000006b3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000832,
      Q => blk00000003_sig00000850
    );
  blk00000003_blk000006b2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000831,
      Q => blk00000003_sig0000084f
    );
  blk00000003_blk000006b1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000830,
      Q => blk00000003_sig0000084e
    );
  blk00000003_blk000006b0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000082f,
      Q => blk00000003_sig0000084d
    );
  blk00000003_blk000006af : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000082e,
      Q => blk00000003_sig0000084c
    );
  blk00000003_blk000006ae : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000082d,
      Q => blk00000003_sig0000084b
    );
  blk00000003_blk000006ad : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000082c,
      Q => blk00000003_sig0000084a
    );
  blk00000003_blk000006ac : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000082b,
      Q => blk00000003_sig00000849
    );
  blk00000003_blk000006ab : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000082a,
      Q => blk00000003_sig00000848
    );
  blk00000003_blk000006aa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000829,
      Q => blk00000003_sig00000847
    );
  blk00000003_blk000006a9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000828,
      Q => blk00000003_sig00000435
    );
  blk00000003_blk000006a8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006aa,
      Q => blk00000003_sig00000846
    );
  blk00000003_blk000006a7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000827,
      Q => blk00000003_sig00000845
    );
  blk00000003_blk000006a6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000826,
      Q => blk00000003_sig00000844
    );
  blk00000003_blk000006a5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000825,
      Q => blk00000003_sig00000843
    );
  blk00000003_blk000006a4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000824,
      Q => blk00000003_sig00000842
    );
  blk00000003_blk000006a3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000823,
      Q => blk00000003_sig00000841
    );
  blk00000003_blk000006a2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000822,
      Q => blk00000003_sig00000840
    );
  blk00000003_blk000006a1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000821,
      Q => blk00000003_sig0000083f
    );
  blk00000003_blk000006a0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000820,
      Q => blk00000003_sig0000083e
    );
  blk00000003_blk0000069f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000081f,
      Q => blk00000003_sig0000083d
    );
  blk00000003_blk0000069e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000081e,
      Q => blk00000003_sig0000083c
    );
  blk00000003_blk0000069d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000081d,
      Q => blk00000003_sig0000083b
    );
  blk00000003_blk0000069c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000081c,
      Q => blk00000003_sig0000083a
    );
  blk00000003_blk0000069b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000081b,
      Q => blk00000003_sig00000839
    );
  blk00000003_blk0000069a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000081a,
      Q => blk00000003_sig00000838
    );
  blk00000003_blk00000699 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000819,
      Q => blk00000003_sig00000837
    );
  blk00000003_blk00000698 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000818,
      Q => blk00000003_sig00000836
    );
  blk00000003_blk00000697 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000817,
      Q => blk00000003_sig00000835
    );
  blk00000003_blk00000696 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000816,
      Q => blk00000003_sig00000834
    );
  blk00000003_blk00000695 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000815,
      Q => blk00000003_sig00000833
    );
  blk00000003_blk00000694 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000814,
      Q => blk00000003_sig00000832
    );
  blk00000003_blk00000693 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000813,
      Q => blk00000003_sig00000831
    );
  blk00000003_blk00000692 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000812,
      Q => blk00000003_sig00000830
    );
  blk00000003_blk00000691 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000811,
      Q => blk00000003_sig0000082f
    );
  blk00000003_blk00000690 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000810,
      Q => blk00000003_sig0000082e
    );
  blk00000003_blk0000068f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000080f,
      Q => blk00000003_sig0000082d
    );
  blk00000003_blk0000068e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000080e,
      Q => blk00000003_sig0000082c
    );
  blk00000003_blk0000068d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000080d,
      Q => blk00000003_sig0000082b
    );
  blk00000003_blk0000068c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000080c,
      Q => blk00000003_sig0000082a
    );
  blk00000003_blk0000068b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000080b,
      Q => blk00000003_sig00000829
    );
  blk00000003_blk0000068a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000080a,
      Q => blk00000003_sig00000828
    );
  blk00000003_blk00000689 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000809,
      Q => blk00000003_sig0000040f
    );
  blk00000003_blk00000688 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ab,
      Q => blk00000003_sig00000827
    );
  blk00000003_blk00000687 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000808,
      Q => blk00000003_sig00000826
    );
  blk00000003_blk00000686 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000807,
      Q => blk00000003_sig00000825
    );
  blk00000003_blk00000685 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000806,
      Q => blk00000003_sig00000824
    );
  blk00000003_blk00000684 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000805,
      Q => blk00000003_sig00000823
    );
  blk00000003_blk00000683 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000804,
      Q => blk00000003_sig00000822
    );
  blk00000003_blk00000682 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000803,
      Q => blk00000003_sig00000821
    );
  blk00000003_blk00000681 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000802,
      Q => blk00000003_sig00000820
    );
  blk00000003_blk00000680 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000801,
      Q => blk00000003_sig0000081f
    );
  blk00000003_blk0000067f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000800,
      Q => blk00000003_sig0000081e
    );
  blk00000003_blk0000067e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007ff,
      Q => blk00000003_sig0000081d
    );
  blk00000003_blk0000067d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007fe,
      Q => blk00000003_sig0000081c
    );
  blk00000003_blk0000067c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007fd,
      Q => blk00000003_sig0000081b
    );
  blk00000003_blk0000067b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007fc,
      Q => blk00000003_sig0000081a
    );
  blk00000003_blk0000067a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007fb,
      Q => blk00000003_sig00000819
    );
  blk00000003_blk00000679 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007fa,
      Q => blk00000003_sig00000818
    );
  blk00000003_blk00000678 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007f9,
      Q => blk00000003_sig00000817
    );
  blk00000003_blk00000677 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007f8,
      Q => blk00000003_sig00000816
    );
  blk00000003_blk00000676 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007f7,
      Q => blk00000003_sig00000815
    );
  blk00000003_blk00000675 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007f6,
      Q => blk00000003_sig00000814
    );
  blk00000003_blk00000674 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007f5,
      Q => blk00000003_sig00000813
    );
  blk00000003_blk00000673 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007f4,
      Q => blk00000003_sig00000812
    );
  blk00000003_blk00000672 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007f3,
      Q => blk00000003_sig00000811
    );
  blk00000003_blk00000671 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007f2,
      Q => blk00000003_sig00000810
    );
  blk00000003_blk00000670 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007f1,
      Q => blk00000003_sig0000080f
    );
  blk00000003_blk0000066f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007f0,
      Q => blk00000003_sig0000080e
    );
  blk00000003_blk0000066e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007ef,
      Q => blk00000003_sig0000080d
    );
  blk00000003_blk0000066d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007ee,
      Q => blk00000003_sig0000080c
    );
  blk00000003_blk0000066c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007ed,
      Q => blk00000003_sig0000080b
    );
  blk00000003_blk0000066b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007ec,
      Q => blk00000003_sig0000080a
    );
  blk00000003_blk0000066a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007eb,
      Q => blk00000003_sig00000809
    );
  blk00000003_blk00000669 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007ea,
      Q => blk00000003_sig000003e9
    );
  blk00000003_blk00000668 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ac,
      Q => blk00000003_sig00000808
    );
  blk00000003_blk00000667 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007e9,
      Q => blk00000003_sig00000807
    );
  blk00000003_blk00000666 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007e8,
      Q => blk00000003_sig00000806
    );
  blk00000003_blk00000665 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007e7,
      Q => blk00000003_sig00000805
    );
  blk00000003_blk00000664 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007e6,
      Q => blk00000003_sig00000804
    );
  blk00000003_blk00000663 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007e5,
      Q => blk00000003_sig00000803
    );
  blk00000003_blk00000662 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007e4,
      Q => blk00000003_sig00000802
    );
  blk00000003_blk00000661 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007e3,
      Q => blk00000003_sig00000801
    );
  blk00000003_blk00000660 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007e2,
      Q => blk00000003_sig00000800
    );
  blk00000003_blk0000065f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007e1,
      Q => blk00000003_sig000007ff
    );
  blk00000003_blk0000065e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007e0,
      Q => blk00000003_sig000007fe
    );
  blk00000003_blk0000065d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007df,
      Q => blk00000003_sig000007fd
    );
  blk00000003_blk0000065c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007de,
      Q => blk00000003_sig000007fc
    );
  blk00000003_blk0000065b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007dd,
      Q => blk00000003_sig000007fb
    );
  blk00000003_blk0000065a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007dc,
      Q => blk00000003_sig000007fa
    );
  blk00000003_blk00000659 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007db,
      Q => blk00000003_sig000007f9
    );
  blk00000003_blk00000658 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007da,
      Q => blk00000003_sig000007f8
    );
  blk00000003_blk00000657 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007d9,
      Q => blk00000003_sig000007f7
    );
  blk00000003_blk00000656 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007d8,
      Q => blk00000003_sig000007f6
    );
  blk00000003_blk00000655 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007d7,
      Q => blk00000003_sig000007f5
    );
  blk00000003_blk00000654 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007d6,
      Q => blk00000003_sig000007f4
    );
  blk00000003_blk00000653 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007d5,
      Q => blk00000003_sig000007f3
    );
  blk00000003_blk00000652 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007d4,
      Q => blk00000003_sig000007f2
    );
  blk00000003_blk00000651 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007d3,
      Q => blk00000003_sig000007f1
    );
  blk00000003_blk00000650 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007d2,
      Q => blk00000003_sig000007f0
    );
  blk00000003_blk0000064f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007d1,
      Q => blk00000003_sig000007ef
    );
  blk00000003_blk0000064e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007d0,
      Q => blk00000003_sig000007ee
    );
  blk00000003_blk0000064d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007cf,
      Q => blk00000003_sig000007ed
    );
  blk00000003_blk0000064c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007ce,
      Q => blk00000003_sig000007ec
    );
  blk00000003_blk0000064b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007cd,
      Q => blk00000003_sig000007eb
    );
  blk00000003_blk0000064a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007cc,
      Q => blk00000003_sig000007ea
    );
  blk00000003_blk00000649 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007cb,
      Q => blk00000003_sig000003c3
    );
  blk00000003_blk00000648 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ad,
      Q => blk00000003_sig000007e9
    );
  blk00000003_blk00000647 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007ca,
      Q => blk00000003_sig000007e8
    );
  blk00000003_blk00000646 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007c9,
      Q => blk00000003_sig000007e7
    );
  blk00000003_blk00000645 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007c8,
      Q => blk00000003_sig000007e6
    );
  blk00000003_blk00000644 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007c7,
      Q => blk00000003_sig000007e5
    );
  blk00000003_blk00000643 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007c6,
      Q => blk00000003_sig000007e4
    );
  blk00000003_blk00000642 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007c5,
      Q => blk00000003_sig000007e3
    );
  blk00000003_blk00000641 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007c4,
      Q => blk00000003_sig000007e2
    );
  blk00000003_blk00000640 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007c3,
      Q => blk00000003_sig000007e1
    );
  blk00000003_blk0000063f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007c2,
      Q => blk00000003_sig000007e0
    );
  blk00000003_blk0000063e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007c1,
      Q => blk00000003_sig000007df
    );
  blk00000003_blk0000063d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007c0,
      Q => blk00000003_sig000007de
    );
  blk00000003_blk0000063c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007bf,
      Q => blk00000003_sig000007dd
    );
  blk00000003_blk0000063b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007be,
      Q => blk00000003_sig000007dc
    );
  blk00000003_blk0000063a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007bd,
      Q => blk00000003_sig000007db
    );
  blk00000003_blk00000639 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007bc,
      Q => blk00000003_sig000007da
    );
  blk00000003_blk00000638 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007bb,
      Q => blk00000003_sig000007d9
    );
  blk00000003_blk00000637 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007ba,
      Q => blk00000003_sig000007d8
    );
  blk00000003_blk00000636 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007b9,
      Q => blk00000003_sig000007d7
    );
  blk00000003_blk00000635 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007b8,
      Q => blk00000003_sig000007d6
    );
  blk00000003_blk00000634 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007b7,
      Q => blk00000003_sig000007d5
    );
  blk00000003_blk00000633 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007b6,
      Q => blk00000003_sig000007d4
    );
  blk00000003_blk00000632 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007b5,
      Q => blk00000003_sig000007d3
    );
  blk00000003_blk00000631 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007b4,
      Q => blk00000003_sig000007d2
    );
  blk00000003_blk00000630 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007b3,
      Q => blk00000003_sig000007d1
    );
  blk00000003_blk0000062f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007b2,
      Q => blk00000003_sig000007d0
    );
  blk00000003_blk0000062e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007b1,
      Q => blk00000003_sig000007cf
    );
  blk00000003_blk0000062d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007b0,
      Q => blk00000003_sig000007ce
    );
  blk00000003_blk0000062c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007af,
      Q => blk00000003_sig000007cd
    );
  blk00000003_blk0000062b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007ae,
      Q => blk00000003_sig000007cc
    );
  blk00000003_blk0000062a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007ad,
      Q => blk00000003_sig000007cb
    );
  blk00000003_blk00000629 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007ac,
      Q => blk00000003_sig0000039d
    );
  blk00000003_blk00000628 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ae,
      Q => blk00000003_sig000007ca
    );
  blk00000003_blk00000627 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006c1,
      Q => blk00000003_sig000007c9
    );
  blk00000003_blk00000626 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006c0,
      Q => blk00000003_sig000007c8
    );
  blk00000003_blk00000625 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006be,
      Q => blk00000003_sig000007c7
    );
  blk00000003_blk00000624 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006bc,
      Q => blk00000003_sig000007c6
    );
  blk00000003_blk00000623 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ba,
      Q => blk00000003_sig000007c5
    );
  blk00000003_blk00000622 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006b8,
      Q => blk00000003_sig000007c4
    );
  blk00000003_blk00000621 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006b6,
      Q => blk00000003_sig000007c3
    );
  blk00000003_blk00000620 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006b4,
      Q => blk00000003_sig000007c2
    );
  blk00000003_blk0000061f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006b2,
      Q => blk00000003_sig000007c1
    );
  blk00000003_blk0000061e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007ab,
      Q => blk00000003_sig000007c0
    );
  blk00000003_blk0000061d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007aa,
      Q => blk00000003_sig000007bf
    );
  blk00000003_blk0000061c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007a9,
      Q => blk00000003_sig000007be
    );
  blk00000003_blk0000061b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007a8,
      Q => blk00000003_sig000007bd
    );
  blk00000003_blk0000061a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007a7,
      Q => blk00000003_sig000007bc
    );
  blk00000003_blk00000619 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007a6,
      Q => blk00000003_sig000007bb
    );
  blk00000003_blk00000618 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007a5,
      Q => blk00000003_sig000007ba
    );
  blk00000003_blk00000617 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007a4,
      Q => blk00000003_sig000007b9
    );
  blk00000003_blk00000616 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007a3,
      Q => blk00000003_sig000007b8
    );
  blk00000003_blk00000615 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007a2,
      Q => blk00000003_sig000007b7
    );
  blk00000003_blk00000614 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007a1,
      Q => blk00000003_sig000007b6
    );
  blk00000003_blk00000613 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007a0,
      Q => blk00000003_sig000007b5
    );
  blk00000003_blk00000612 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000079f,
      Q => blk00000003_sig000007b4
    );
  blk00000003_blk00000611 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000079e,
      Q => blk00000003_sig000007b3
    );
  blk00000003_blk00000610 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000079d,
      Q => blk00000003_sig000007b2
    );
  blk00000003_blk0000060f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000079c,
      Q => blk00000003_sig000007b1
    );
  blk00000003_blk0000060e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000079b,
      Q => blk00000003_sig000007b0
    );
  blk00000003_blk0000060d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000079a,
      Q => blk00000003_sig000007af
    );
  blk00000003_blk0000060c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000799,
      Q => blk00000003_sig000007ae
    );
  blk00000003_blk0000060b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000798,
      Q => blk00000003_sig000007ad
    );
  blk00000003_blk0000060a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000797,
      Q => blk00000003_sig000007ac
    );
  blk00000003_blk00000609 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000796,
      Q => blk00000003_sig00000377
    );
  blk00000003_blk00000608 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000795,
      Q => blk00000003_sig000007ab
    );
  blk00000003_blk00000607 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000794,
      Q => blk00000003_sig000007aa
    );
  blk00000003_blk00000606 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000793,
      Q => blk00000003_sig000007a9
    );
  blk00000003_blk00000605 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000792,
      Q => blk00000003_sig000007a8
    );
  blk00000003_blk00000604 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000791,
      Q => blk00000003_sig000007a7
    );
  blk00000003_blk00000603 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000790,
      Q => blk00000003_sig000007a6
    );
  blk00000003_blk00000602 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000078f,
      Q => blk00000003_sig000007a5
    );
  blk00000003_blk00000601 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000078e,
      Q => blk00000003_sig000007a4
    );
  blk00000003_blk00000600 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000078d,
      Q => blk00000003_sig000007a3
    );
  blk00000003_blk000005ff : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000078c,
      Q => blk00000003_sig000007a2
    );
  blk00000003_blk000005fe : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000078b,
      Q => blk00000003_sig000007a1
    );
  blk00000003_blk000005fd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000078a,
      Q => blk00000003_sig000007a0
    );
  blk00000003_blk000005fc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000789,
      Q => blk00000003_sig0000079f
    );
  blk00000003_blk000005fb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000788,
      Q => blk00000003_sig0000079e
    );
  blk00000003_blk000005fa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000787,
      Q => blk00000003_sig0000079d
    );
  blk00000003_blk000005f9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000786,
      Q => blk00000003_sig0000079c
    );
  blk00000003_blk000005f8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000785,
      Q => blk00000003_sig0000079b
    );
  blk00000003_blk000005f7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000784,
      Q => blk00000003_sig0000079a
    );
  blk00000003_blk000005f6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000783,
      Q => blk00000003_sig00000799
    );
  blk00000003_blk000005f5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000782,
      Q => blk00000003_sig00000798
    );
  blk00000003_blk000005f4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000781,
      Q => blk00000003_sig00000797
    );
  blk00000003_blk000005f3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000780,
      Q => blk00000003_sig00000796
    );
  blk00000003_blk000005f2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000077f,
      Q => blk00000003_sig00000351
    );
  blk00000003_blk000005f1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006b0,
      Q => blk00000003_sig000006bf
    );
  blk00000003_blk000005f0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000078,
      Q => blk00000003_sig000006bd
    );
  blk00000003_blk000005ef : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007a,
      Q => blk00000003_sig000006bb
    );
  blk00000003_blk000005ee : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007c,
      Q => blk00000003_sig000006b9
    );
  blk00000003_blk000005ed : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007e,
      Q => blk00000003_sig000006b7
    );
  blk00000003_blk000005ec : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000080,
      Q => blk00000003_sig000006b5
    );
  blk00000003_blk000005eb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000082,
      Q => blk00000003_sig000006b3
    );
  blk00000003_blk000005ea : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000084,
      Q => blk00000003_sig000006b1
    );
  blk00000003_blk000005e9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000077e,
      Q => blk00000003_sig00000795
    );
  blk00000003_blk000005e8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000077d,
      Q => blk00000003_sig00000794
    );
  blk00000003_blk000005e7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000077c,
      Q => blk00000003_sig00000793
    );
  blk00000003_blk000005e6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000077b,
      Q => blk00000003_sig00000792
    );
  blk00000003_blk000005e5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000077a,
      Q => blk00000003_sig00000791
    );
  blk00000003_blk000005e4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000779,
      Q => blk00000003_sig00000790
    );
  blk00000003_blk000005e3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000778,
      Q => blk00000003_sig0000078f
    );
  blk00000003_blk000005e2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000777,
      Q => blk00000003_sig0000078e
    );
  blk00000003_blk000005e1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000776,
      Q => blk00000003_sig0000078d
    );
  blk00000003_blk000005e0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000775,
      Q => blk00000003_sig0000078c
    );
  blk00000003_blk000005df : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000774,
      Q => blk00000003_sig0000078b
    );
  blk00000003_blk000005de : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000773,
      Q => blk00000003_sig0000078a
    );
  blk00000003_blk000005dd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000772,
      Q => blk00000003_sig00000789
    );
  blk00000003_blk000005dc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000771,
      Q => blk00000003_sig00000788
    );
  blk00000003_blk000005db : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000770,
      Q => blk00000003_sig00000787
    );
  blk00000003_blk000005da : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000076f,
      Q => blk00000003_sig00000786
    );
  blk00000003_blk000005d9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000076e,
      Q => blk00000003_sig00000785
    );
  blk00000003_blk000005d8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000076d,
      Q => blk00000003_sig00000784
    );
  blk00000003_blk000005d7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000076c,
      Q => blk00000003_sig00000783
    );
  blk00000003_blk000005d6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000076b,
      Q => blk00000003_sig00000782
    );
  blk00000003_blk000005d5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000076a,
      Q => blk00000003_sig00000781
    );
  blk00000003_blk000005d4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000769,
      Q => blk00000003_sig00000780
    );
  blk00000003_blk000005d3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000768,
      Q => blk00000003_sig0000077f
    );
  blk00000003_blk000005d2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000767,
      Q => blk00000003_sig0000032b
    );
  blk00000003_blk000005d1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000766,
      Q => blk00000003_sig0000077e
    );
  blk00000003_blk000005d0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000765,
      Q => blk00000003_sig0000077d
    );
  blk00000003_blk000005cf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000764,
      Q => blk00000003_sig0000077c
    );
  blk00000003_blk000005ce : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000763,
      Q => blk00000003_sig0000077b
    );
  blk00000003_blk000005cd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000762,
      Q => blk00000003_sig0000077a
    );
  blk00000003_blk000005cc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000761,
      Q => blk00000003_sig00000779
    );
  blk00000003_blk000005cb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000760,
      Q => blk00000003_sig00000778
    );
  blk00000003_blk000005ca : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000075f,
      Q => blk00000003_sig00000777
    );
  blk00000003_blk000005c9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000075e,
      Q => blk00000003_sig00000776
    );
  blk00000003_blk000005c8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000075d,
      Q => blk00000003_sig00000775
    );
  blk00000003_blk000005c7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000075c,
      Q => blk00000003_sig00000774
    );
  blk00000003_blk000005c6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000075b,
      Q => blk00000003_sig00000773
    );
  blk00000003_blk000005c5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000075a,
      Q => blk00000003_sig00000772
    );
  blk00000003_blk000005c4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000759,
      Q => blk00000003_sig00000771
    );
  blk00000003_blk000005c3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000758,
      Q => blk00000003_sig00000770
    );
  blk00000003_blk000005c2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000757,
      Q => blk00000003_sig0000076f
    );
  blk00000003_blk000005c1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000756,
      Q => blk00000003_sig0000076e
    );
  blk00000003_blk000005c0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000755,
      Q => blk00000003_sig0000076d
    );
  blk00000003_blk000005bf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000754,
      Q => blk00000003_sig0000076c
    );
  blk00000003_blk000005be : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000753,
      Q => blk00000003_sig0000076b
    );
  blk00000003_blk000005bd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000752,
      Q => blk00000003_sig0000076a
    );
  blk00000003_blk000005bc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000751,
      Q => blk00000003_sig00000769
    );
  blk00000003_blk000005bb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000750,
      Q => blk00000003_sig00000768
    );
  blk00000003_blk000005ba : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000074f,
      Q => blk00000003_sig00000767
    );
  blk00000003_blk000005b9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000074e,
      Q => blk00000003_sig00000305
    );
  blk00000003_blk000005b8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000074d,
      Q => blk00000003_sig00000766
    );
  blk00000003_blk000005b7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000074c,
      Q => blk00000003_sig00000765
    );
  blk00000003_blk000005b6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000074b,
      Q => blk00000003_sig00000764
    );
  blk00000003_blk000005b5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000074a,
      Q => blk00000003_sig00000763
    );
  blk00000003_blk000005b4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000749,
      Q => blk00000003_sig00000762
    );
  blk00000003_blk000005b3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000748,
      Q => blk00000003_sig00000761
    );
  blk00000003_blk000005b2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000747,
      Q => blk00000003_sig00000760
    );
  blk00000003_blk000005b1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000746,
      Q => blk00000003_sig0000075f
    );
  blk00000003_blk000005b0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000745,
      Q => blk00000003_sig0000075e
    );
  blk00000003_blk000005af : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000744,
      Q => blk00000003_sig0000075d
    );
  blk00000003_blk000005ae : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000743,
      Q => blk00000003_sig0000075c
    );
  blk00000003_blk000005ad : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000742,
      Q => blk00000003_sig0000075b
    );
  blk00000003_blk000005ac : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000741,
      Q => blk00000003_sig0000075a
    );
  blk00000003_blk000005ab : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000740,
      Q => blk00000003_sig00000759
    );
  blk00000003_blk000005aa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000073f,
      Q => blk00000003_sig00000758
    );
  blk00000003_blk000005a9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000073e,
      Q => blk00000003_sig00000757
    );
  blk00000003_blk000005a8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000073d,
      Q => blk00000003_sig00000756
    );
  blk00000003_blk000005a7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000073c,
      Q => blk00000003_sig00000755
    );
  blk00000003_blk000005a6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000073b,
      Q => blk00000003_sig00000754
    );
  blk00000003_blk000005a5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000073a,
      Q => blk00000003_sig00000753
    );
  blk00000003_blk000005a4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000739,
      Q => blk00000003_sig00000752
    );
  blk00000003_blk000005a3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000738,
      Q => blk00000003_sig00000751
    );
  blk00000003_blk000005a2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000737,
      Q => blk00000003_sig00000750
    );
  blk00000003_blk000005a1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000736,
      Q => blk00000003_sig0000074f
    );
  blk00000003_blk000005a0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000735,
      Q => blk00000003_sig0000074e
    );
  blk00000003_blk0000059f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000734,
      Q => blk00000003_sig000002df
    );
  blk00000003_blk0000059e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000733,
      Q => blk00000003_sig0000074d
    );
  blk00000003_blk0000059d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000732,
      Q => blk00000003_sig0000074c
    );
  blk00000003_blk0000059c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000731,
      Q => blk00000003_sig0000074b
    );
  blk00000003_blk0000059b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000730,
      Q => blk00000003_sig0000074a
    );
  blk00000003_blk0000059a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000072f,
      Q => blk00000003_sig00000749
    );
  blk00000003_blk00000599 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000072e,
      Q => blk00000003_sig00000748
    );
  blk00000003_blk00000598 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000072d,
      Q => blk00000003_sig00000747
    );
  blk00000003_blk00000597 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000072c,
      Q => blk00000003_sig00000746
    );
  blk00000003_blk00000596 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000072b,
      Q => blk00000003_sig00000745
    );
  blk00000003_blk00000595 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000072a,
      Q => blk00000003_sig00000744
    );
  blk00000003_blk00000594 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000729,
      Q => blk00000003_sig00000743
    );
  blk00000003_blk00000593 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000728,
      Q => blk00000003_sig00000742
    );
  blk00000003_blk00000592 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000727,
      Q => blk00000003_sig00000741
    );
  blk00000003_blk00000591 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000726,
      Q => blk00000003_sig00000740
    );
  blk00000003_blk00000590 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000725,
      Q => blk00000003_sig0000073f
    );
  blk00000003_blk0000058f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000724,
      Q => blk00000003_sig0000073e
    );
  blk00000003_blk0000058e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000723,
      Q => blk00000003_sig0000073d
    );
  blk00000003_blk0000058d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000722,
      Q => blk00000003_sig0000073c
    );
  blk00000003_blk0000058c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000721,
      Q => blk00000003_sig0000073b
    );
  blk00000003_blk0000058b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000720,
      Q => blk00000003_sig0000073a
    );
  blk00000003_blk0000058a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000071f,
      Q => blk00000003_sig00000739
    );
  blk00000003_blk00000589 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000071e,
      Q => blk00000003_sig00000738
    );
  blk00000003_blk00000588 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000071d,
      Q => blk00000003_sig00000737
    );
  blk00000003_blk00000587 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000071c,
      Q => blk00000003_sig00000736
    );
  blk00000003_blk00000586 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000071b,
      Q => blk00000003_sig00000735
    );
  blk00000003_blk00000585 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000071a,
      Q => blk00000003_sig00000734
    );
  blk00000003_blk00000584 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000719,
      Q => blk00000003_sig000002b9
    );
  blk00000003_blk00000583 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000718,
      Q => blk00000003_sig00000733
    );
  blk00000003_blk00000582 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000717,
      Q => blk00000003_sig00000732
    );
  blk00000003_blk00000581 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000716,
      Q => blk00000003_sig00000731
    );
  blk00000003_blk00000580 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000715,
      Q => blk00000003_sig00000730
    );
  blk00000003_blk0000057f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000714,
      Q => blk00000003_sig0000072f
    );
  blk00000003_blk0000057e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000713,
      Q => blk00000003_sig0000072e
    );
  blk00000003_blk0000057d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000712,
      Q => blk00000003_sig0000072d
    );
  blk00000003_blk0000057c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000711,
      Q => blk00000003_sig0000072c
    );
  blk00000003_blk0000057b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000710,
      Q => blk00000003_sig0000072b
    );
  blk00000003_blk0000057a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000070f,
      Q => blk00000003_sig0000072a
    );
  blk00000003_blk00000579 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000070e,
      Q => blk00000003_sig00000729
    );
  blk00000003_blk00000578 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000070d,
      Q => blk00000003_sig00000728
    );
  blk00000003_blk00000577 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000070c,
      Q => blk00000003_sig00000727
    );
  blk00000003_blk00000576 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000070b,
      Q => blk00000003_sig00000726
    );
  blk00000003_blk00000575 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000070a,
      Q => blk00000003_sig00000725
    );
  blk00000003_blk00000574 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000709,
      Q => blk00000003_sig00000724
    );
  blk00000003_blk00000573 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000708,
      Q => blk00000003_sig00000723
    );
  blk00000003_blk00000572 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000707,
      Q => blk00000003_sig00000722
    );
  blk00000003_blk00000571 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000706,
      Q => blk00000003_sig00000721
    );
  blk00000003_blk00000570 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000705,
      Q => blk00000003_sig00000720
    );
  blk00000003_blk0000056f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000704,
      Q => blk00000003_sig0000071f
    );
  blk00000003_blk0000056e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000703,
      Q => blk00000003_sig0000071e
    );
  blk00000003_blk0000056d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000702,
      Q => blk00000003_sig0000071d
    );
  blk00000003_blk0000056c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000701,
      Q => blk00000003_sig0000071c
    );
  blk00000003_blk0000056b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000700,
      Q => blk00000003_sig0000071b
    );
  blk00000003_blk0000056a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ff,
      Q => blk00000003_sig0000071a
    );
  blk00000003_blk00000569 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006fe,
      Q => blk00000003_sig00000719
    );
  blk00000003_blk00000568 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006fd,
      Q => blk00000003_sig00000293
    );
  blk00000003_blk00000567 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006fc,
      Q => blk00000003_sig00000718
    );
  blk00000003_blk00000566 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006fb,
      Q => blk00000003_sig00000717
    );
  blk00000003_blk00000565 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006fa,
      Q => blk00000003_sig00000716
    );
  blk00000003_blk00000564 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006f9,
      Q => blk00000003_sig00000715
    );
  blk00000003_blk00000563 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006f8,
      Q => blk00000003_sig00000714
    );
  blk00000003_blk00000562 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006f7,
      Q => blk00000003_sig00000713
    );
  blk00000003_blk00000561 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006f6,
      Q => blk00000003_sig00000712
    );
  blk00000003_blk00000560 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006f5,
      Q => blk00000003_sig00000711
    );
  blk00000003_blk0000055f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006f4,
      Q => blk00000003_sig00000710
    );
  blk00000003_blk0000055e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006f3,
      Q => blk00000003_sig0000070f
    );
  blk00000003_blk0000055d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006f2,
      Q => blk00000003_sig0000070e
    );
  blk00000003_blk0000055c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006f1,
      Q => blk00000003_sig0000070d
    );
  blk00000003_blk0000055b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006f0,
      Q => blk00000003_sig0000070c
    );
  blk00000003_blk0000055a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ef,
      Q => blk00000003_sig0000070b
    );
  blk00000003_blk00000559 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ee,
      Q => blk00000003_sig0000070a
    );
  blk00000003_blk00000558 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ed,
      Q => blk00000003_sig00000709
    );
  blk00000003_blk00000557 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ec,
      Q => blk00000003_sig00000708
    );
  blk00000003_blk00000556 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006eb,
      Q => blk00000003_sig00000707
    );
  blk00000003_blk00000555 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ea,
      Q => blk00000003_sig00000706
    );
  blk00000003_blk00000554 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006e9,
      Q => blk00000003_sig00000705
    );
  blk00000003_blk00000553 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006e8,
      Q => blk00000003_sig00000704
    );
  blk00000003_blk00000552 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006e7,
      Q => blk00000003_sig00000703
    );
  blk00000003_blk00000551 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006e6,
      Q => blk00000003_sig00000702
    );
  blk00000003_blk00000550 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006e5,
      Q => blk00000003_sig00000701
    );
  blk00000003_blk0000054f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006e4,
      Q => blk00000003_sig00000700
    );
  blk00000003_blk0000054e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006e3,
      Q => blk00000003_sig000006ff
    );
  blk00000003_blk0000054d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006e2,
      Q => blk00000003_sig000006fe
    );
  blk00000003_blk0000054c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006e1,
      Q => blk00000003_sig000006fd
    );
  blk00000003_blk0000054b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006e0,
      Q => blk00000003_sig0000026d
    );
  blk00000003_blk0000054a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006df,
      Q => blk00000003_sig000006fc
    );
  blk00000003_blk00000549 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006de,
      Q => blk00000003_sig000006fb
    );
  blk00000003_blk00000548 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006dd,
      Q => blk00000003_sig000006fa
    );
  blk00000003_blk00000547 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006dc,
      Q => blk00000003_sig000006f9
    );
  blk00000003_blk00000546 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006db,
      Q => blk00000003_sig000006f8
    );
  blk00000003_blk00000545 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006da,
      Q => blk00000003_sig000006f7
    );
  blk00000003_blk00000544 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006d9,
      Q => blk00000003_sig000006f6
    );
  blk00000003_blk00000543 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006d8,
      Q => blk00000003_sig000006f5
    );
  blk00000003_blk00000542 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006d7,
      Q => blk00000003_sig000006f4
    );
  blk00000003_blk00000541 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006d6,
      Q => blk00000003_sig000006f3
    );
  blk00000003_blk00000540 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006d5,
      Q => blk00000003_sig000006f2
    );
  blk00000003_blk0000053f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006d4,
      Q => blk00000003_sig000006f1
    );
  blk00000003_blk0000053e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006d3,
      Q => blk00000003_sig000006f0
    );
  blk00000003_blk0000053d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006d2,
      Q => blk00000003_sig000006ef
    );
  blk00000003_blk0000053c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006d1,
      Q => blk00000003_sig000006ee
    );
  blk00000003_blk0000053b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006d0,
      Q => blk00000003_sig000006ed
    );
  blk00000003_blk0000053a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006cf,
      Q => blk00000003_sig000006ec
    );
  blk00000003_blk00000539 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ce,
      Q => blk00000003_sig000006eb
    );
  blk00000003_blk00000538 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006cd,
      Q => blk00000003_sig000006ea
    );
  blk00000003_blk00000537 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006cc,
      Q => blk00000003_sig000006e9
    );
  blk00000003_blk00000536 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006cb,
      Q => blk00000003_sig000006e8
    );
  blk00000003_blk00000535 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ca,
      Q => blk00000003_sig000006e7
    );
  blk00000003_blk00000534 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006c9,
      Q => blk00000003_sig000006e6
    );
  blk00000003_blk00000533 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006c8,
      Q => blk00000003_sig000006e5
    );
  blk00000003_blk00000532 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006c7,
      Q => blk00000003_sig000006e4
    );
  blk00000003_blk00000531 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006c6,
      Q => blk00000003_sig000006e3
    );
  blk00000003_blk00000530 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006c5,
      Q => blk00000003_sig000006e2
    );
  blk00000003_blk0000052f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006c4,
      Q => blk00000003_sig000006e1
    );
  blk00000003_blk0000052e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006c3,
      Q => blk00000003_sig000006e0
    );
  blk00000003_blk0000052d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006c2,
      Q => blk00000003_sig00000247
    );
  blk00000003_blk0000052c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000da,
      Q => blk00000003_sig000006df
    );
  blk00000003_blk0000052b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d9,
      Q => blk00000003_sig000006de
    );
  blk00000003_blk0000052a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d8,
      Q => blk00000003_sig000006dd
    );
  blk00000003_blk00000529 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d7,
      Q => blk00000003_sig000006dc
    );
  blk00000003_blk00000528 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d6,
      Q => blk00000003_sig000006db
    );
  blk00000003_blk00000527 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d5,
      Q => blk00000003_sig000006da
    );
  blk00000003_blk00000526 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d4,
      Q => blk00000003_sig000006d9
    );
  blk00000003_blk00000525 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d3,
      Q => blk00000003_sig000006d8
    );
  blk00000003_blk00000524 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d2,
      Q => blk00000003_sig000006d7
    );
  blk00000003_blk00000523 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d1,
      Q => blk00000003_sig000006d6
    );
  blk00000003_blk00000522 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d0,
      Q => blk00000003_sig000006d5
    );
  blk00000003_blk00000521 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000cf,
      Q => blk00000003_sig000006d4
    );
  blk00000003_blk00000520 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ce,
      Q => blk00000003_sig000006d3
    );
  blk00000003_blk0000051f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000cd,
      Q => blk00000003_sig000006d2
    );
  blk00000003_blk0000051e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000cc,
      Q => blk00000003_sig000006d1
    );
  blk00000003_blk0000051d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000cb,
      Q => blk00000003_sig000006d0
    );
  blk00000003_blk0000051c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ca,
      Q => blk00000003_sig000006cf
    );
  blk00000003_blk0000051b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c9,
      Q => blk00000003_sig000006ce
    );
  blk00000003_blk0000051a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c8,
      Q => blk00000003_sig000006cd
    );
  blk00000003_blk00000519 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c7,
      Q => blk00000003_sig000006cc
    );
  blk00000003_blk00000518 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c6,
      Q => blk00000003_sig000006cb
    );
  blk00000003_blk00000517 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c5,
      Q => blk00000003_sig000006ca
    );
  blk00000003_blk00000516 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c4,
      Q => blk00000003_sig000006c9
    );
  blk00000003_blk00000515 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c3,
      Q => blk00000003_sig000006c8
    );
  blk00000003_blk00000514 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c2,
      Q => blk00000003_sig000006c7
    );
  blk00000003_blk00000513 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c1,
      Q => blk00000003_sig000006c6
    );
  blk00000003_blk00000512 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c0,
      Q => blk00000003_sig000006c5
    );
  blk00000003_blk00000511 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000bf,
      Q => blk00000003_sig000006c4
    );
  blk00000003_blk00000510 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000be,
      Q => blk00000003_sig000006c3
    );
  blk00000003_blk0000050f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000bd,
      Q => blk00000003_sig000006c2
    );
  blk00000003_blk0000050e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000bc,
      Q => blk00000003_sig00000221
    );
  blk00000003_blk0000050d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006af,
      Q => blk00000003_sig000006c1
    );
  blk00000003_blk0000050c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006bf,
      Q => blk00000003_sig000006c0
    );
  blk00000003_blk0000050b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006bd,
      Q => blk00000003_sig000006be
    );
  blk00000003_blk0000050a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006bb,
      Q => blk00000003_sig000006bc
    );
  blk00000003_blk00000509 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006b9,
      Q => blk00000003_sig000006ba
    );
  blk00000003_blk00000508 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006b7,
      Q => blk00000003_sig000006b8
    );
  blk00000003_blk00000507 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006b5,
      Q => blk00000003_sig000006b6
    );
  blk00000003_blk00000506 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006b3,
      Q => blk00000003_sig000006b4
    );
  blk00000003_blk00000505 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006b1,
      Q => blk00000003_sig000006b2
    );
  blk00000003_blk00000504 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001fb,
      Q => blk00000003_sig0000021b
    );
  blk00000003_blk00000503 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001f8,
      Q => blk00000003_sig0000021a
    );
  blk00000003_blk00000502 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001f5,
      Q => blk00000003_sig00000219
    );
  blk00000003_blk00000501 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001f2,
      Q => blk00000003_sig00000218
    );
  blk00000003_blk00000500 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001ef,
      Q => blk00000003_sig00000217
    );
  blk00000003_blk000004ff : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001ec,
      Q => blk00000003_sig00000216
    );
  blk00000003_blk000004fe : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001e9,
      Q => blk00000003_sig00000215
    );
  blk00000003_blk000004fd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001e6,
      Q => blk00000003_sig0000021c
    );
  blk00000003_blk000004fc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000220,
      Q => blk00000003_sig00000241
    );
  blk00000003_blk000004fb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000214,
      Q => blk00000003_sig00000240
    );
  blk00000003_blk000004fa : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000211,
      Q => blk00000003_sig0000023f
    );
  blk00000003_blk000004f9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000020e,
      Q => blk00000003_sig0000023e
    );
  blk00000003_blk000004f8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000020b,
      Q => blk00000003_sig0000023d
    );
  blk00000003_blk000004f7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000208,
      Q => blk00000003_sig0000023c
    );
  blk00000003_blk000004f6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000205,
      Q => blk00000003_sig0000023b
    );
  blk00000003_blk000004f5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000202,
      Q => blk00000003_sig00000242
    );
  blk00000003_blk000004f4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001ff,
      Q => blk00000003_sig00000097
    );
  blk00000003_blk000004f3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000246,
      Q => blk00000003_sig00000267
    );
  blk00000003_blk000004f2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000023a,
      Q => blk00000003_sig00000266
    );
  blk00000003_blk000004f1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000237,
      Q => blk00000003_sig00000265
    );
  blk00000003_blk000004f0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000234,
      Q => blk00000003_sig00000264
    );
  blk00000003_blk000004ef : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000231,
      Q => blk00000003_sig00000263
    );
  blk00000003_blk000004ee : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000022e,
      Q => blk00000003_sig00000262
    );
  blk00000003_blk000004ed : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000022b,
      Q => blk00000003_sig00000261
    );
  blk00000003_blk000004ec : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000228,
      Q => blk00000003_sig00000268
    );
  blk00000003_blk000004eb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000225,
      Q => blk00000003_sig00000094
    );
  blk00000003_blk000004ea : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000026c,
      Q => blk00000003_sig0000028d
    );
  blk00000003_blk000004e9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000260,
      Q => blk00000003_sig0000028c
    );
  blk00000003_blk000004e8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000025d,
      Q => blk00000003_sig0000028b
    );
  blk00000003_blk000004e7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000025a,
      Q => blk00000003_sig0000028a
    );
  blk00000003_blk000004e6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000257,
      Q => blk00000003_sig00000289
    );
  blk00000003_blk000004e5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000254,
      Q => blk00000003_sig00000288
    );
  blk00000003_blk000004e4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000251,
      Q => blk00000003_sig00000287
    );
  blk00000003_blk000004e3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000024e,
      Q => blk00000003_sig0000028e
    );
  blk00000003_blk000004e2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000024b,
      Q => blk00000003_sig00000090
    );
  blk00000003_blk000004e1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000292,
      Q => blk00000003_sig000002b3
    );
  blk00000003_blk000004e0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000286,
      Q => blk00000003_sig000002b2
    );
  blk00000003_blk000004df : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000283,
      Q => blk00000003_sig000002b1
    );
  blk00000003_blk000004de : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000280,
      Q => blk00000003_sig000002b0
    );
  blk00000003_blk000004dd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000027d,
      Q => blk00000003_sig000002af
    );
  blk00000003_blk000004dc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000027a,
      Q => blk00000003_sig000002ae
    );
  blk00000003_blk000004db : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000277,
      Q => blk00000003_sig000002ad
    );
  blk00000003_blk000004da : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000274,
      Q => blk00000003_sig000002b4
    );
  blk00000003_blk000004d9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000271,
      Q => blk00000003_sig0000008b
    );
  blk00000003_blk000004d8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002b8,
      Q => blk00000003_sig000002d9
    );
  blk00000003_blk000004d7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002ac,
      Q => blk00000003_sig000002d8
    );
  blk00000003_blk000004d6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002a9,
      Q => blk00000003_sig000002d7
    );
  blk00000003_blk000004d5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002a6,
      Q => blk00000003_sig000002d6
    );
  blk00000003_blk000004d4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002a3,
      Q => blk00000003_sig000002d5
    );
  blk00000003_blk000004d3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002a0,
      Q => blk00000003_sig000002d4
    );
  blk00000003_blk000004d2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000029d,
      Q => blk00000003_sig000002d3
    );
  blk00000003_blk000004d1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000029a,
      Q => blk00000003_sig000002da
    );
  blk00000003_blk000004d0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000297,
      Q => blk00000003_sig00000085
    );
  blk00000003_blk000004cf : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002de,
      Q => blk00000003_sig000002ff
    );
  blk00000003_blk000004ce : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002d2,
      Q => blk00000003_sig000002fe
    );
  blk00000003_blk000004cd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002cf,
      Q => blk00000003_sig000002fd
    );
  blk00000003_blk000004cc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002cc,
      Q => blk00000003_sig000002fc
    );
  blk00000003_blk000004cb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002c9,
      Q => blk00000003_sig000002fb
    );
  blk00000003_blk000004ca : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002c6,
      Q => blk00000003_sig000002fa
    );
  blk00000003_blk000004c9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002c3,
      Q => blk00000003_sig000002f9
    );
  blk00000003_blk000004c8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002c0,
      Q => blk00000003_sig00000300
    );
  blk00000003_blk000004c7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002bd,
      Q => blk00000003_sig00000077
    );
  blk00000003_blk000004c6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000304,
      Q => blk00000003_sig00000325
    );
  blk00000003_blk000004c5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002f8,
      Q => blk00000003_sig00000324
    );
  blk00000003_blk000004c4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002f5,
      Q => blk00000003_sig00000323
    );
  blk00000003_blk000004c3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002f2,
      Q => blk00000003_sig00000322
    );
  blk00000003_blk000004c2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002ef,
      Q => blk00000003_sig00000321
    );
  blk00000003_blk000004c1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002ec,
      Q => blk00000003_sig00000320
    );
  blk00000003_blk000004c0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002e9,
      Q => blk00000003_sig0000031f
    );
  blk00000003_blk000004bf : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002e6,
      Q => blk00000003_sig00000326
    );
  blk00000003_blk000004be : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002e3,
      Q => blk00000003_sig000006b0
    );
  blk00000003_blk000004bd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000032a,
      Q => blk00000003_sig0000034b
    );
  blk00000003_blk000004bc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000031e,
      Q => blk00000003_sig0000034a
    );
  blk00000003_blk000004bb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000031b,
      Q => blk00000003_sig00000349
    );
  blk00000003_blk000004ba : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000318,
      Q => blk00000003_sig00000348
    );
  blk00000003_blk000004b9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000315,
      Q => blk00000003_sig00000347
    );
  blk00000003_blk000004b8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000312,
      Q => blk00000003_sig00000346
    );
  blk00000003_blk000004b7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000030f,
      Q => blk00000003_sig00000345
    );
  blk00000003_blk000004b6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000030c,
      Q => blk00000003_sig0000034c
    );
  blk00000003_blk000004b5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000309,
      Q => blk00000003_sig000006af
    );
  blk00000003_blk000004b4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000350,
      Q => blk00000003_sig00000371
    );
  blk00000003_blk000004b3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000344,
      Q => blk00000003_sig00000370
    );
  blk00000003_blk000004b2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000341,
      Q => blk00000003_sig0000036f
    );
  blk00000003_blk000004b1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000033e,
      Q => blk00000003_sig0000036e
    );
  blk00000003_blk000004b0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000033b,
      Q => blk00000003_sig0000036d
    );
  blk00000003_blk000004af : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000338,
      Q => blk00000003_sig0000036c
    );
  blk00000003_blk000004ae : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000335,
      Q => blk00000003_sig0000036b
    );
  blk00000003_blk000004ad : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000332,
      Q => blk00000003_sig00000372
    );
  blk00000003_blk000004ac : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000032f,
      Q => blk00000003_sig000006ae
    );
  blk00000003_blk000004ab : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000376,
      Q => blk00000003_sig00000397
    );
  blk00000003_blk000004aa : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000036a,
      Q => blk00000003_sig00000396
    );
  blk00000003_blk000004a9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000367,
      Q => blk00000003_sig00000395
    );
  blk00000003_blk000004a8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000364,
      Q => blk00000003_sig00000394
    );
  blk00000003_blk000004a7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000361,
      Q => blk00000003_sig00000393
    );
  blk00000003_blk000004a6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000035e,
      Q => blk00000003_sig00000392
    );
  blk00000003_blk000004a5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000035b,
      Q => blk00000003_sig00000391
    );
  blk00000003_blk000004a4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000358,
      Q => blk00000003_sig00000398
    );
  blk00000003_blk000004a3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000355,
      Q => blk00000003_sig000006ad
    );
  blk00000003_blk000004a2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000039c,
      Q => blk00000003_sig000003bd
    );
  blk00000003_blk000004a1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000390,
      Q => blk00000003_sig000003bc
    );
  blk00000003_blk000004a0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000038d,
      Q => blk00000003_sig000003bb
    );
  blk00000003_blk0000049f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000038a,
      Q => blk00000003_sig000003ba
    );
  blk00000003_blk0000049e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000387,
      Q => blk00000003_sig000003b9
    );
  blk00000003_blk0000049d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000384,
      Q => blk00000003_sig000003b8
    );
  blk00000003_blk0000049c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000381,
      Q => blk00000003_sig000003b7
    );
  blk00000003_blk0000049b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000037e,
      Q => blk00000003_sig000003be
    );
  blk00000003_blk0000049a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000037b,
      Q => blk00000003_sig000006ac
    );
  blk00000003_blk00000499 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003c2,
      Q => blk00000003_sig000003e3
    );
  blk00000003_blk00000498 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003b6,
      Q => blk00000003_sig000003e2
    );
  blk00000003_blk00000497 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003b3,
      Q => blk00000003_sig000003e1
    );
  blk00000003_blk00000496 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003b0,
      Q => blk00000003_sig000003e0
    );
  blk00000003_blk00000495 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003ad,
      Q => blk00000003_sig000003df
    );
  blk00000003_blk00000494 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003aa,
      Q => blk00000003_sig000003de
    );
  blk00000003_blk00000493 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003a7,
      Q => blk00000003_sig000003dd
    );
  blk00000003_blk00000492 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003a4,
      Q => blk00000003_sig000003e4
    );
  blk00000003_blk00000491 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003a1,
      Q => blk00000003_sig000006ab
    );
  blk00000003_blk00000490 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003e8,
      Q => blk00000003_sig00000409
    );
  blk00000003_blk0000048f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003dc,
      Q => blk00000003_sig00000408
    );
  blk00000003_blk0000048e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003d9,
      Q => blk00000003_sig00000407
    );
  blk00000003_blk0000048d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003d6,
      Q => blk00000003_sig00000406
    );
  blk00000003_blk0000048c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003d3,
      Q => blk00000003_sig00000405
    );
  blk00000003_blk0000048b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003d0,
      Q => blk00000003_sig00000404
    );
  blk00000003_blk0000048a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003cd,
      Q => blk00000003_sig00000403
    );
  blk00000003_blk00000489 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003ca,
      Q => blk00000003_sig0000040a
    );
  blk00000003_blk00000488 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003c7,
      Q => blk00000003_sig000006aa
    );
  blk00000003_blk00000487 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000040e,
      Q => blk00000003_sig0000042f
    );
  blk00000003_blk00000486 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000402,
      Q => blk00000003_sig0000042e
    );
  blk00000003_blk00000485 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003ff,
      Q => blk00000003_sig0000042d
    );
  blk00000003_blk00000484 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003fc,
      Q => blk00000003_sig0000042c
    );
  blk00000003_blk00000483 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003f9,
      Q => blk00000003_sig0000042b
    );
  blk00000003_blk00000482 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003f6,
      Q => blk00000003_sig0000042a
    );
  blk00000003_blk00000481 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003f3,
      Q => blk00000003_sig00000429
    );
  blk00000003_blk00000480 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003f0,
      Q => blk00000003_sig00000430
    );
  blk00000003_blk0000047f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003ed,
      Q => blk00000003_sig000006a9
    );
  blk00000003_blk0000047e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000434,
      Q => blk00000003_sig00000455
    );
  blk00000003_blk0000047d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000428,
      Q => blk00000003_sig00000454
    );
  blk00000003_blk0000047c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000425,
      Q => blk00000003_sig00000453
    );
  blk00000003_blk0000047b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000422,
      Q => blk00000003_sig00000452
    );
  blk00000003_blk0000047a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000041f,
      Q => blk00000003_sig00000451
    );
  blk00000003_blk00000479 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000041c,
      Q => blk00000003_sig00000450
    );
  blk00000003_blk00000478 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000419,
      Q => blk00000003_sig0000044f
    );
  blk00000003_blk00000477 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000416,
      Q => blk00000003_sig00000456
    );
  blk00000003_blk00000476 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000413,
      Q => blk00000003_sig000006a8
    );
  blk00000003_blk00000475 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000045a,
      Q => blk00000003_sig0000047b
    );
  blk00000003_blk00000474 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000044e,
      Q => blk00000003_sig0000047a
    );
  blk00000003_blk00000473 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000044b,
      Q => blk00000003_sig00000479
    );
  blk00000003_blk00000472 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000448,
      Q => blk00000003_sig00000478
    );
  blk00000003_blk00000471 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000445,
      Q => blk00000003_sig00000477
    );
  blk00000003_blk00000470 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000442,
      Q => blk00000003_sig00000476
    );
  blk00000003_blk0000046f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000043f,
      Q => blk00000003_sig00000475
    );
  blk00000003_blk0000046e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000043c,
      Q => blk00000003_sig0000047c
    );
  blk00000003_blk0000046d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000439,
      Q => blk00000003_sig000006a7
    );
  blk00000003_blk0000046c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000480,
      Q => blk00000003_sig000004a1
    );
  blk00000003_blk0000046b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000474,
      Q => blk00000003_sig000004a0
    );
  blk00000003_blk0000046a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000471,
      Q => blk00000003_sig0000049f
    );
  blk00000003_blk00000469 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000046e,
      Q => blk00000003_sig0000049e
    );
  blk00000003_blk00000468 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000046b,
      Q => blk00000003_sig0000049d
    );
  blk00000003_blk00000467 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000468,
      Q => blk00000003_sig0000049c
    );
  blk00000003_blk00000466 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000465,
      Q => blk00000003_sig0000049b
    );
  blk00000003_blk00000465 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000462,
      Q => blk00000003_sig000004a2
    );
  blk00000003_blk00000464 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000045f,
      Q => blk00000003_sig000006a6
    );
  blk00000003_blk00000463 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004a6,
      Q => blk00000003_sig000004c7
    );
  blk00000003_blk00000462 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000049a,
      Q => blk00000003_sig000004c6
    );
  blk00000003_blk00000461 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000497,
      Q => blk00000003_sig000004c5
    );
  blk00000003_blk00000460 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000494,
      Q => blk00000003_sig000004c4
    );
  blk00000003_blk0000045f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000491,
      Q => blk00000003_sig000004c3
    );
  blk00000003_blk0000045e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000048e,
      Q => blk00000003_sig000004c2
    );
  blk00000003_blk0000045d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000048b,
      Q => blk00000003_sig000004c1
    );
  blk00000003_blk0000045c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000488,
      Q => blk00000003_sig000004c8
    );
  blk00000003_blk0000045b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000485,
      Q => blk00000003_sig000006a5
    );
  blk00000003_blk0000045a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004cc,
      Q => blk00000003_sig000004ed
    );
  blk00000003_blk00000459 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004c0,
      Q => blk00000003_sig000004ec
    );
  blk00000003_blk00000458 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004bd,
      Q => blk00000003_sig000004eb
    );
  blk00000003_blk00000457 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004ba,
      Q => blk00000003_sig000004ea
    );
  blk00000003_blk00000456 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004b7,
      Q => blk00000003_sig000004e9
    );
  blk00000003_blk00000455 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004b4,
      Q => blk00000003_sig000004e8
    );
  blk00000003_blk00000454 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004b1,
      Q => blk00000003_sig000004e7
    );
  blk00000003_blk00000453 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004ae,
      Q => blk00000003_sig000004ee
    );
  blk00000003_blk00000452 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004ab,
      Q => blk00000003_sig000006a4
    );
  blk00000003_blk00000451 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004f2,
      Q => blk00000003_sig00000513
    );
  blk00000003_blk00000450 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004e6,
      Q => blk00000003_sig00000512
    );
  blk00000003_blk0000044f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004e3,
      Q => blk00000003_sig00000511
    );
  blk00000003_blk0000044e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004e0,
      Q => blk00000003_sig00000510
    );
  blk00000003_blk0000044d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004dd,
      Q => blk00000003_sig0000050f
    );
  blk00000003_blk0000044c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004da,
      Q => blk00000003_sig0000050e
    );
  blk00000003_blk0000044b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004d7,
      Q => blk00000003_sig0000050d
    );
  blk00000003_blk0000044a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004d4,
      Q => blk00000003_sig00000514
    );
  blk00000003_blk00000449 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004d1,
      Q => blk00000003_sig000006a3
    );
  blk00000003_blk00000448 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000518,
      Q => blk00000003_sig00000539
    );
  blk00000003_blk00000447 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000050c,
      Q => blk00000003_sig00000538
    );
  blk00000003_blk00000446 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000509,
      Q => blk00000003_sig00000537
    );
  blk00000003_blk00000445 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000506,
      Q => blk00000003_sig00000536
    );
  blk00000003_blk00000444 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000503,
      Q => blk00000003_sig00000535
    );
  blk00000003_blk00000443 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000500,
      Q => blk00000003_sig00000534
    );
  blk00000003_blk00000442 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004fd,
      Q => blk00000003_sig00000533
    );
  blk00000003_blk00000441 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004fa,
      Q => blk00000003_sig0000053a
    );
  blk00000003_blk00000440 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004f7,
      Q => blk00000003_sig000006a2
    );
  blk00000003_blk0000043f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000053e,
      Q => blk00000003_sig0000055f
    );
  blk00000003_blk0000043e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000532,
      Q => blk00000003_sig0000055e
    );
  blk00000003_blk0000043d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000052f,
      Q => blk00000003_sig0000055d
    );
  blk00000003_blk0000043c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000052c,
      Q => blk00000003_sig0000055c
    );
  blk00000003_blk0000043b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000529,
      Q => blk00000003_sig0000055b
    );
  blk00000003_blk0000043a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000526,
      Q => blk00000003_sig0000055a
    );
  blk00000003_blk00000439 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000523,
      Q => blk00000003_sig00000559
    );
  blk00000003_blk00000438 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000520,
      Q => blk00000003_sig00000560
    );
  blk00000003_blk00000437 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000051d,
      Q => blk00000003_sig000006a1
    );
  blk00000003_blk00000436 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000564,
      Q => blk00000003_sig00000585
    );
  blk00000003_blk00000435 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000558,
      Q => blk00000003_sig00000584
    );
  blk00000003_blk00000434 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000555,
      Q => blk00000003_sig00000583
    );
  blk00000003_blk00000433 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000552,
      Q => blk00000003_sig00000582
    );
  blk00000003_blk00000432 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000054f,
      Q => blk00000003_sig00000581
    );
  blk00000003_blk00000431 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000054c,
      Q => blk00000003_sig00000580
    );
  blk00000003_blk00000430 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000549,
      Q => blk00000003_sig0000057f
    );
  blk00000003_blk0000042f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000546,
      Q => blk00000003_sig00000586
    );
  blk00000003_blk0000042e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000543,
      Q => blk00000003_sig000006a0
    );
  blk00000003_blk0000042d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000058a,
      Q => blk00000003_sig000005ab
    );
  blk00000003_blk0000042c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000057e,
      Q => blk00000003_sig000005aa
    );
  blk00000003_blk0000042b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000057b,
      Q => blk00000003_sig000005a9
    );
  blk00000003_blk0000042a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000578,
      Q => blk00000003_sig000005a8
    );
  blk00000003_blk00000429 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000575,
      Q => blk00000003_sig000005a7
    );
  blk00000003_blk00000428 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000572,
      Q => blk00000003_sig000005a6
    );
  blk00000003_blk00000427 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000056f,
      Q => blk00000003_sig000005a5
    );
  blk00000003_blk00000426 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000056c,
      Q => blk00000003_sig000005ac
    );
  blk00000003_blk00000425 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000569,
      Q => blk00000003_sig0000069f
    );
  blk00000003_blk00000424 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005b0,
      Q => blk00000003_sig000005d0
    );
  blk00000003_blk00000423 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005a4,
      Q => blk00000003_sig000005cf
    );
  blk00000003_blk00000422 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005a1,
      Q => blk00000003_sig000005ce
    );
  blk00000003_blk00000421 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000059e,
      Q => blk00000003_sig000005cd
    );
  blk00000003_blk00000420 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000059b,
      Q => blk00000003_sig000005cc
    );
  blk00000003_blk0000041f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000598,
      Q => blk00000003_sig000005cb
    );
  blk00000003_blk0000041e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000595,
      Q => blk00000003_sig000005ca
    );
  blk00000003_blk0000041d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000592,
      Q => blk00000003_sig000005d1
    );
  blk00000003_blk0000041c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000058f,
      Q => blk00000003_sig0000069e
    );
  blk00000003_blk0000041b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005d5,
      Q => blk00000003_sig000005f5
    );
  blk00000003_blk0000041a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005c9,
      Q => blk00000003_sig000005f4
    );
  blk00000003_blk00000419 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005c6,
      Q => blk00000003_sig000005f3
    );
  blk00000003_blk00000418 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005c3,
      Q => blk00000003_sig000005f2
    );
  blk00000003_blk00000417 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005c0,
      Q => blk00000003_sig000005f1
    );
  blk00000003_blk00000416 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005bd,
      Q => blk00000003_sig000005f0
    );
  blk00000003_blk00000415 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005ba,
      Q => blk00000003_sig000005ef
    );
  blk00000003_blk00000414 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005b7,
      Q => blk00000003_sig000005f6
    );
  blk00000003_blk00000413 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005b4,
      Q => blk00000003_sig0000069d
    );
  blk00000003_blk00000412 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005fa,
      Q => blk00000003_sig0000061a
    );
  blk00000003_blk00000411 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005ee,
      Q => blk00000003_sig00000619
    );
  blk00000003_blk00000410 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005eb,
      Q => blk00000003_sig00000618
    );
  blk00000003_blk0000040f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005e8,
      Q => blk00000003_sig00000617
    );
  blk00000003_blk0000040e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005e5,
      Q => blk00000003_sig00000616
    );
  blk00000003_blk0000040d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005e2,
      Q => blk00000003_sig00000615
    );
  blk00000003_blk0000040c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005df,
      Q => blk00000003_sig00000614
    );
  blk00000003_blk0000040b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005dc,
      Q => blk00000003_sig0000061b
    );
  blk00000003_blk0000040a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005d9,
      Q => blk00000003_sig0000069c
    );
  blk00000003_blk00000409 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000061f,
      Q => blk00000003_sig0000063f
    );
  blk00000003_blk00000408 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000613,
      Q => blk00000003_sig0000063e
    );
  blk00000003_blk00000407 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000610,
      Q => blk00000003_sig0000063d
    );
  blk00000003_blk00000406 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000060d,
      Q => blk00000003_sig0000063c
    );
  blk00000003_blk00000405 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000060a,
      Q => blk00000003_sig0000063b
    );
  blk00000003_blk00000404 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000607,
      Q => blk00000003_sig0000063a
    );
  blk00000003_blk00000403 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000604,
      Q => blk00000003_sig00000639
    );
  blk00000003_blk00000402 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000601,
      Q => blk00000003_sig00000640
    );
  blk00000003_blk00000401 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005fe,
      Q => blk00000003_sig0000069b
    );
  blk00000003_blk00000400 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000644,
      Q => blk00000003_sig00000664
    );
  blk00000003_blk000003ff : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000638,
      Q => blk00000003_sig00000663
    );
  blk00000003_blk000003fe : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000635,
      Q => blk00000003_sig00000662
    );
  blk00000003_blk000003fd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000632,
      Q => blk00000003_sig00000661
    );
  blk00000003_blk000003fc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000062f,
      Q => blk00000003_sig00000660
    );
  blk00000003_blk000003fb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000062c,
      Q => blk00000003_sig0000065f
    );
  blk00000003_blk000003fa : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000629,
      Q => blk00000003_sig0000065e
    );
  blk00000003_blk000003f9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000626,
      Q => blk00000003_sig00000665
    );
  blk00000003_blk000003f8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000623,
      Q => blk00000003_sig0000069a
    );
  blk00000003_blk000003f7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000669,
      Q => blk00000003_sig00000689
    );
  blk00000003_blk000003f6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000065d,
      Q => blk00000003_sig00000688
    );
  blk00000003_blk000003f5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000065a,
      Q => blk00000003_sig00000687
    );
  blk00000003_blk000003f4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000657,
      Q => blk00000003_sig00000686
    );
  blk00000003_blk000003f3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000654,
      Q => blk00000003_sig00000685
    );
  blk00000003_blk000003f2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000651,
      Q => blk00000003_sig00000684
    );
  blk00000003_blk000003f1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000064e,
      Q => blk00000003_sig00000683
    );
  blk00000003_blk000003f0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000064b,
      Q => blk00000003_sig0000068a
    );
  blk00000003_blk000003ef : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000648,
      Q => blk00000003_sig00000699
    );
  blk00000003_blk000003ee : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000068e,
      Q => blk00000003_sig00000698
    );
  blk00000003_blk000003ed : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000682,
      Q => blk00000003_sig00000697
    );
  blk00000003_blk000003ec : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000067f,
      Q => blk00000003_sig00000696
    );
  blk00000003_blk000003eb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000067c,
      Q => blk00000003_sig00000695
    );
  blk00000003_blk000003ea : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000679,
      Q => blk00000003_sig00000694
    );
  blk00000003_blk000003e9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000676,
      Q => blk00000003_sig00000693
    );
  blk00000003_blk000003e8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000673,
      Q => blk00000003_sig00000692
    );
  blk00000003_blk000003e7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000670,
      Q => blk00000003_sig00000691
    );
  blk00000003_blk000003e6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000066d,
      Q => blk00000003_sig00000690
    );
  blk00000003_blk000003e5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000068b,
      Q => blk00000003_sig0000068f
    );
  blk00000003_blk000003e4 : MUXCY
    port map (
      CI => blk00000003_sig0000068c,
      DI => blk00000003_sig0000009a,
      S => blk00000003_sig0000068d,
      O => blk00000003_sig00000680
    );
  blk00000003_blk000003e3 : XORCY
    port map (
      CI => blk00000003_sig0000068c,
      LI => blk00000003_sig0000068d,
      O => blk00000003_sig0000068e
    );
  blk00000003_blk000003e2 : MUXCY
    port map (
      CI => blk00000003_sig0000066b,
      DI => blk00000003_sig0000068a,
      S => blk00000003_sig0000066c,
      O => blk00000003_sig0000068b
    );
  blk00000003_blk000003e1 : MUXCY
    port map (
      CI => blk00000003_sig00000680,
      DI => blk00000003_sig00000689,
      S => blk00000003_sig00000681,
      O => blk00000003_sig0000067d
    );
  blk00000003_blk000003e0 : MUXCY
    port map (
      CI => blk00000003_sig0000067d,
      DI => blk00000003_sig00000688,
      S => blk00000003_sig0000067e,
      O => blk00000003_sig0000067a
    );
  blk00000003_blk000003df : MUXCY
    port map (
      CI => blk00000003_sig0000067a,
      DI => blk00000003_sig00000687,
      S => blk00000003_sig0000067b,
      O => blk00000003_sig00000677
    );
  blk00000003_blk000003de : MUXCY
    port map (
      CI => blk00000003_sig00000677,
      DI => blk00000003_sig00000686,
      S => blk00000003_sig00000678,
      O => blk00000003_sig00000674
    );
  blk00000003_blk000003dd : MUXCY
    port map (
      CI => blk00000003_sig00000674,
      DI => blk00000003_sig00000685,
      S => blk00000003_sig00000675,
      O => blk00000003_sig00000671
    );
  blk00000003_blk000003dc : MUXCY
    port map (
      CI => blk00000003_sig00000671,
      DI => blk00000003_sig00000684,
      S => blk00000003_sig00000672,
      O => blk00000003_sig0000066e
    );
  blk00000003_blk000003db : MUXCY
    port map (
      CI => blk00000003_sig0000066e,
      DI => blk00000003_sig00000683,
      S => blk00000003_sig0000066f,
      O => blk00000003_sig0000066b
    );
  blk00000003_blk000003da : XORCY
    port map (
      CI => blk00000003_sig00000680,
      LI => blk00000003_sig00000681,
      O => blk00000003_sig00000682
    );
  blk00000003_blk000003d9 : XORCY
    port map (
      CI => blk00000003_sig0000067d,
      LI => blk00000003_sig0000067e,
      O => blk00000003_sig0000067f
    );
  blk00000003_blk000003d8 : XORCY
    port map (
      CI => blk00000003_sig0000067a,
      LI => blk00000003_sig0000067b,
      O => blk00000003_sig0000067c
    );
  blk00000003_blk000003d7 : XORCY
    port map (
      CI => blk00000003_sig00000677,
      LI => blk00000003_sig00000678,
      O => blk00000003_sig00000679
    );
  blk00000003_blk000003d6 : XORCY
    port map (
      CI => blk00000003_sig00000674,
      LI => blk00000003_sig00000675,
      O => blk00000003_sig00000676
    );
  blk00000003_blk000003d5 : XORCY
    port map (
      CI => blk00000003_sig00000671,
      LI => blk00000003_sig00000672,
      O => blk00000003_sig00000673
    );
  blk00000003_blk000003d4 : XORCY
    port map (
      CI => blk00000003_sig0000066e,
      LI => blk00000003_sig0000066f,
      O => blk00000003_sig00000670
    );
  blk00000003_blk000003d3 : XORCY
    port map (
      CI => blk00000003_sig0000066b,
      LI => blk00000003_sig0000066c,
      O => blk00000003_sig0000066d
    );
  blk00000003_blk000003d2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000666,
      Q => blk00000003_sig0000066a
    );
  blk00000003_blk000003d1 : MUXCY
    port map (
      CI => blk00000003_sig00000667,
      DI => blk00000003_sig00000058,
      S => blk00000003_sig00000668,
      O => blk00000003_sig0000065b
    );
  blk00000003_blk000003d0 : XORCY
    port map (
      CI => blk00000003_sig00000667,
      LI => blk00000003_sig00000668,
      O => blk00000003_sig00000669
    );
  blk00000003_blk000003cf : MUXCY
    port map (
      CI => blk00000003_sig00000646,
      DI => blk00000003_sig00000665,
      S => blk00000003_sig00000647,
      O => blk00000003_sig00000666
    );
  blk00000003_blk000003ce : MUXCY
    port map (
      CI => blk00000003_sig0000065b,
      DI => blk00000003_sig00000664,
      S => blk00000003_sig0000065c,
      O => blk00000003_sig00000658
    );
  blk00000003_blk000003cd : MUXCY
    port map (
      CI => blk00000003_sig00000658,
      DI => blk00000003_sig00000663,
      S => blk00000003_sig00000659,
      O => blk00000003_sig00000655
    );
  blk00000003_blk000003cc : MUXCY
    port map (
      CI => blk00000003_sig00000655,
      DI => blk00000003_sig00000662,
      S => blk00000003_sig00000656,
      O => blk00000003_sig00000652
    );
  blk00000003_blk000003cb : MUXCY
    port map (
      CI => blk00000003_sig00000652,
      DI => blk00000003_sig00000661,
      S => blk00000003_sig00000653,
      O => blk00000003_sig0000064f
    );
  blk00000003_blk000003ca : MUXCY
    port map (
      CI => blk00000003_sig0000064f,
      DI => blk00000003_sig00000660,
      S => blk00000003_sig00000650,
      O => blk00000003_sig0000064c
    );
  blk00000003_blk000003c9 : MUXCY
    port map (
      CI => blk00000003_sig0000064c,
      DI => blk00000003_sig0000065f,
      S => blk00000003_sig0000064d,
      O => blk00000003_sig00000649
    );
  blk00000003_blk000003c8 : MUXCY
    port map (
      CI => blk00000003_sig00000649,
      DI => blk00000003_sig0000065e,
      S => blk00000003_sig0000064a,
      O => blk00000003_sig00000646
    );
  blk00000003_blk000003c7 : XORCY
    port map (
      CI => blk00000003_sig0000065b,
      LI => blk00000003_sig0000065c,
      O => blk00000003_sig0000065d
    );
  blk00000003_blk000003c6 : XORCY
    port map (
      CI => blk00000003_sig00000658,
      LI => blk00000003_sig00000659,
      O => blk00000003_sig0000065a
    );
  blk00000003_blk000003c5 : XORCY
    port map (
      CI => blk00000003_sig00000655,
      LI => blk00000003_sig00000656,
      O => blk00000003_sig00000657
    );
  blk00000003_blk000003c4 : XORCY
    port map (
      CI => blk00000003_sig00000652,
      LI => blk00000003_sig00000653,
      O => blk00000003_sig00000654
    );
  blk00000003_blk000003c3 : XORCY
    port map (
      CI => blk00000003_sig0000064f,
      LI => blk00000003_sig00000650,
      O => blk00000003_sig00000651
    );
  blk00000003_blk000003c2 : XORCY
    port map (
      CI => blk00000003_sig0000064c,
      LI => blk00000003_sig0000064d,
      O => blk00000003_sig0000064e
    );
  blk00000003_blk000003c1 : XORCY
    port map (
      CI => blk00000003_sig00000649,
      LI => blk00000003_sig0000064a,
      O => blk00000003_sig0000064b
    );
  blk00000003_blk000003c0 : XORCY
    port map (
      CI => blk00000003_sig00000646,
      LI => blk00000003_sig00000647,
      O => blk00000003_sig00000648
    );
  blk00000003_blk000003bf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000641,
      Q => blk00000003_sig00000645
    );
  blk00000003_blk000003be : MUXCY
    port map (
      CI => blk00000003_sig00000642,
      DI => blk00000003_sig0000005c,
      S => blk00000003_sig00000643,
      O => blk00000003_sig00000636
    );
  blk00000003_blk000003bd : XORCY
    port map (
      CI => blk00000003_sig00000642,
      LI => blk00000003_sig00000643,
      O => blk00000003_sig00000644
    );
  blk00000003_blk000003bc : MUXCY
    port map (
      CI => blk00000003_sig00000621,
      DI => blk00000003_sig00000640,
      S => blk00000003_sig00000622,
      O => blk00000003_sig00000641
    );
  blk00000003_blk000003bb : MUXCY
    port map (
      CI => blk00000003_sig00000636,
      DI => blk00000003_sig0000063f,
      S => blk00000003_sig00000637,
      O => blk00000003_sig00000633
    );
  blk00000003_blk000003ba : MUXCY
    port map (
      CI => blk00000003_sig00000633,
      DI => blk00000003_sig0000063e,
      S => blk00000003_sig00000634,
      O => blk00000003_sig00000630
    );
  blk00000003_blk000003b9 : MUXCY
    port map (
      CI => blk00000003_sig00000630,
      DI => blk00000003_sig0000063d,
      S => blk00000003_sig00000631,
      O => blk00000003_sig0000062d
    );
  blk00000003_blk000003b8 : MUXCY
    port map (
      CI => blk00000003_sig0000062d,
      DI => blk00000003_sig0000063c,
      S => blk00000003_sig0000062e,
      O => blk00000003_sig0000062a
    );
  blk00000003_blk000003b7 : MUXCY
    port map (
      CI => blk00000003_sig0000062a,
      DI => blk00000003_sig0000063b,
      S => blk00000003_sig0000062b,
      O => blk00000003_sig00000627
    );
  blk00000003_blk000003b6 : MUXCY
    port map (
      CI => blk00000003_sig00000627,
      DI => blk00000003_sig0000063a,
      S => blk00000003_sig00000628,
      O => blk00000003_sig00000624
    );
  blk00000003_blk000003b5 : MUXCY
    port map (
      CI => blk00000003_sig00000624,
      DI => blk00000003_sig00000639,
      S => blk00000003_sig00000625,
      O => blk00000003_sig00000621
    );
  blk00000003_blk000003b4 : XORCY
    port map (
      CI => blk00000003_sig00000636,
      LI => blk00000003_sig00000637,
      O => blk00000003_sig00000638
    );
  blk00000003_blk000003b3 : XORCY
    port map (
      CI => blk00000003_sig00000633,
      LI => blk00000003_sig00000634,
      O => blk00000003_sig00000635
    );
  blk00000003_blk000003b2 : XORCY
    port map (
      CI => blk00000003_sig00000630,
      LI => blk00000003_sig00000631,
      O => blk00000003_sig00000632
    );
  blk00000003_blk000003b1 : XORCY
    port map (
      CI => blk00000003_sig0000062d,
      LI => blk00000003_sig0000062e,
      O => blk00000003_sig0000062f
    );
  blk00000003_blk000003b0 : XORCY
    port map (
      CI => blk00000003_sig0000062a,
      LI => blk00000003_sig0000062b,
      O => blk00000003_sig0000062c
    );
  blk00000003_blk000003af : XORCY
    port map (
      CI => blk00000003_sig00000627,
      LI => blk00000003_sig00000628,
      O => blk00000003_sig00000629
    );
  blk00000003_blk000003ae : XORCY
    port map (
      CI => blk00000003_sig00000624,
      LI => blk00000003_sig00000625,
      O => blk00000003_sig00000626
    );
  blk00000003_blk000003ad : XORCY
    port map (
      CI => blk00000003_sig00000621,
      LI => blk00000003_sig00000622,
      O => blk00000003_sig00000623
    );
  blk00000003_blk000003ac : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000061c,
      Q => blk00000003_sig00000620
    );
  blk00000003_blk000003ab : MUXCY
    port map (
      CI => blk00000003_sig0000061d,
      DI => blk00000003_sig00000061,
      S => blk00000003_sig0000061e,
      O => blk00000003_sig00000611
    );
  blk00000003_blk000003aa : XORCY
    port map (
      CI => blk00000003_sig0000061d,
      LI => blk00000003_sig0000061e,
      O => blk00000003_sig0000061f
    );
  blk00000003_blk000003a9 : MUXCY
    port map (
      CI => blk00000003_sig000005fc,
      DI => blk00000003_sig0000061b,
      S => blk00000003_sig000005fd,
      O => blk00000003_sig0000061c
    );
  blk00000003_blk000003a8 : MUXCY
    port map (
      CI => blk00000003_sig00000611,
      DI => blk00000003_sig0000061a,
      S => blk00000003_sig00000612,
      O => blk00000003_sig0000060e
    );
  blk00000003_blk000003a7 : MUXCY
    port map (
      CI => blk00000003_sig0000060e,
      DI => blk00000003_sig00000619,
      S => blk00000003_sig0000060f,
      O => blk00000003_sig0000060b
    );
  blk00000003_blk000003a6 : MUXCY
    port map (
      CI => blk00000003_sig0000060b,
      DI => blk00000003_sig00000618,
      S => blk00000003_sig0000060c,
      O => blk00000003_sig00000608
    );
  blk00000003_blk000003a5 : MUXCY
    port map (
      CI => blk00000003_sig00000608,
      DI => blk00000003_sig00000617,
      S => blk00000003_sig00000609,
      O => blk00000003_sig00000605
    );
  blk00000003_blk000003a4 : MUXCY
    port map (
      CI => blk00000003_sig00000605,
      DI => blk00000003_sig00000616,
      S => blk00000003_sig00000606,
      O => blk00000003_sig00000602
    );
  blk00000003_blk000003a3 : MUXCY
    port map (
      CI => blk00000003_sig00000602,
      DI => blk00000003_sig00000615,
      S => blk00000003_sig00000603,
      O => blk00000003_sig000005ff
    );
  blk00000003_blk000003a2 : MUXCY
    port map (
      CI => blk00000003_sig000005ff,
      DI => blk00000003_sig00000614,
      S => blk00000003_sig00000600,
      O => blk00000003_sig000005fc
    );
  blk00000003_blk000003a1 : XORCY
    port map (
      CI => blk00000003_sig00000611,
      LI => blk00000003_sig00000612,
      O => blk00000003_sig00000613
    );
  blk00000003_blk000003a0 : XORCY
    port map (
      CI => blk00000003_sig0000060e,
      LI => blk00000003_sig0000060f,
      O => blk00000003_sig00000610
    );
  blk00000003_blk0000039f : XORCY
    port map (
      CI => blk00000003_sig0000060b,
      LI => blk00000003_sig0000060c,
      O => blk00000003_sig0000060d
    );
  blk00000003_blk0000039e : XORCY
    port map (
      CI => blk00000003_sig00000608,
      LI => blk00000003_sig00000609,
      O => blk00000003_sig0000060a
    );
  blk00000003_blk0000039d : XORCY
    port map (
      CI => blk00000003_sig00000605,
      LI => blk00000003_sig00000606,
      O => blk00000003_sig00000607
    );
  blk00000003_blk0000039c : XORCY
    port map (
      CI => blk00000003_sig00000602,
      LI => blk00000003_sig00000603,
      O => blk00000003_sig00000604
    );
  blk00000003_blk0000039b : XORCY
    port map (
      CI => blk00000003_sig000005ff,
      LI => blk00000003_sig00000600,
      O => blk00000003_sig00000601
    );
  blk00000003_blk0000039a : XORCY
    port map (
      CI => blk00000003_sig000005fc,
      LI => blk00000003_sig000005fd,
      O => blk00000003_sig000005fe
    );
  blk00000003_blk00000399 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005f7,
      Q => blk00000003_sig000005fb
    );
  blk00000003_blk00000398 : MUXCY
    port map (
      CI => blk00000003_sig000005f8,
      DI => blk00000003_sig00000067,
      S => blk00000003_sig000005f9,
      O => blk00000003_sig000005ec
    );
  blk00000003_blk00000397 : XORCY
    port map (
      CI => blk00000003_sig000005f8,
      LI => blk00000003_sig000005f9,
      O => blk00000003_sig000005fa
    );
  blk00000003_blk00000396 : MUXCY
    port map (
      CI => blk00000003_sig000005d7,
      DI => blk00000003_sig000005f6,
      S => blk00000003_sig000005d8,
      O => blk00000003_sig000005f7
    );
  blk00000003_blk00000395 : MUXCY
    port map (
      CI => blk00000003_sig000005ec,
      DI => blk00000003_sig000005f5,
      S => blk00000003_sig000005ed,
      O => blk00000003_sig000005e9
    );
  blk00000003_blk00000394 : MUXCY
    port map (
      CI => blk00000003_sig000005e9,
      DI => blk00000003_sig000005f4,
      S => blk00000003_sig000005ea,
      O => blk00000003_sig000005e6
    );
  blk00000003_blk00000393 : MUXCY
    port map (
      CI => blk00000003_sig000005e6,
      DI => blk00000003_sig000005f3,
      S => blk00000003_sig000005e7,
      O => blk00000003_sig000005e3
    );
  blk00000003_blk00000392 : MUXCY
    port map (
      CI => blk00000003_sig000005e3,
      DI => blk00000003_sig000005f2,
      S => blk00000003_sig000005e4,
      O => blk00000003_sig000005e0
    );
  blk00000003_blk00000391 : MUXCY
    port map (
      CI => blk00000003_sig000005e0,
      DI => blk00000003_sig000005f1,
      S => blk00000003_sig000005e1,
      O => blk00000003_sig000005dd
    );
  blk00000003_blk00000390 : MUXCY
    port map (
      CI => blk00000003_sig000005dd,
      DI => blk00000003_sig000005f0,
      S => blk00000003_sig000005de,
      O => blk00000003_sig000005da
    );
  blk00000003_blk0000038f : MUXCY
    port map (
      CI => blk00000003_sig000005da,
      DI => blk00000003_sig000005ef,
      S => blk00000003_sig000005db,
      O => blk00000003_sig000005d7
    );
  blk00000003_blk0000038e : XORCY
    port map (
      CI => blk00000003_sig000005ec,
      LI => blk00000003_sig000005ed,
      O => blk00000003_sig000005ee
    );
  blk00000003_blk0000038d : XORCY
    port map (
      CI => blk00000003_sig000005e9,
      LI => blk00000003_sig000005ea,
      O => blk00000003_sig000005eb
    );
  blk00000003_blk0000038c : XORCY
    port map (
      CI => blk00000003_sig000005e6,
      LI => blk00000003_sig000005e7,
      O => blk00000003_sig000005e8
    );
  blk00000003_blk0000038b : XORCY
    port map (
      CI => blk00000003_sig000005e3,
      LI => blk00000003_sig000005e4,
      O => blk00000003_sig000005e5
    );
  blk00000003_blk0000038a : XORCY
    port map (
      CI => blk00000003_sig000005e0,
      LI => blk00000003_sig000005e1,
      O => blk00000003_sig000005e2
    );
  blk00000003_blk00000389 : XORCY
    port map (
      CI => blk00000003_sig000005dd,
      LI => blk00000003_sig000005de,
      O => blk00000003_sig000005df
    );
  blk00000003_blk00000388 : XORCY
    port map (
      CI => blk00000003_sig000005da,
      LI => blk00000003_sig000005db,
      O => blk00000003_sig000005dc
    );
  blk00000003_blk00000387 : XORCY
    port map (
      CI => blk00000003_sig000005d7,
      LI => blk00000003_sig000005d8,
      O => blk00000003_sig000005d9
    );
  blk00000003_blk00000386 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005d2,
      Q => blk00000003_sig000005d6
    );
  blk00000003_blk00000385 : MUXCY
    port map (
      CI => blk00000003_sig000005d3,
      DI => blk00000003_sig0000006e,
      S => blk00000003_sig000005d4,
      O => blk00000003_sig000005c7
    );
  blk00000003_blk00000384 : XORCY
    port map (
      CI => blk00000003_sig000005d3,
      LI => blk00000003_sig000005d4,
      O => blk00000003_sig000005d5
    );
  blk00000003_blk00000383 : MUXCY
    port map (
      CI => blk00000003_sig000005b2,
      DI => blk00000003_sig000005d1,
      S => blk00000003_sig000005b3,
      O => blk00000003_sig000005d2
    );
  blk00000003_blk00000382 : MUXCY
    port map (
      CI => blk00000003_sig000005c7,
      DI => blk00000003_sig000005d0,
      S => blk00000003_sig000005c8,
      O => blk00000003_sig000005c4
    );
  blk00000003_blk00000381 : MUXCY
    port map (
      CI => blk00000003_sig000005c4,
      DI => blk00000003_sig000005cf,
      S => blk00000003_sig000005c5,
      O => blk00000003_sig000005c1
    );
  blk00000003_blk00000380 : MUXCY
    port map (
      CI => blk00000003_sig000005c1,
      DI => blk00000003_sig000005ce,
      S => blk00000003_sig000005c2,
      O => blk00000003_sig000005be
    );
  blk00000003_blk0000037f : MUXCY
    port map (
      CI => blk00000003_sig000005be,
      DI => blk00000003_sig000005cd,
      S => blk00000003_sig000005bf,
      O => blk00000003_sig000005bb
    );
  blk00000003_blk0000037e : MUXCY
    port map (
      CI => blk00000003_sig000005bb,
      DI => blk00000003_sig000005cc,
      S => blk00000003_sig000005bc,
      O => blk00000003_sig000005b8
    );
  blk00000003_blk0000037d : MUXCY
    port map (
      CI => blk00000003_sig000005b8,
      DI => blk00000003_sig000005cb,
      S => blk00000003_sig000005b9,
      O => blk00000003_sig000005b5
    );
  blk00000003_blk0000037c : MUXCY
    port map (
      CI => blk00000003_sig000005b5,
      DI => blk00000003_sig000005ca,
      S => blk00000003_sig000005b6,
      O => blk00000003_sig000005b2
    );
  blk00000003_blk0000037b : XORCY
    port map (
      CI => blk00000003_sig000005c7,
      LI => blk00000003_sig000005c8,
      O => blk00000003_sig000005c9
    );
  blk00000003_blk0000037a : XORCY
    port map (
      CI => blk00000003_sig000005c4,
      LI => blk00000003_sig000005c5,
      O => blk00000003_sig000005c6
    );
  blk00000003_blk00000379 : XORCY
    port map (
      CI => blk00000003_sig000005c1,
      LI => blk00000003_sig000005c2,
      O => blk00000003_sig000005c3
    );
  blk00000003_blk00000378 : XORCY
    port map (
      CI => blk00000003_sig000005be,
      LI => blk00000003_sig000005bf,
      O => blk00000003_sig000005c0
    );
  blk00000003_blk00000377 : XORCY
    port map (
      CI => blk00000003_sig000005bb,
      LI => blk00000003_sig000005bc,
      O => blk00000003_sig000005bd
    );
  blk00000003_blk00000376 : XORCY
    port map (
      CI => blk00000003_sig000005b8,
      LI => blk00000003_sig000005b9,
      O => blk00000003_sig000005ba
    );
  blk00000003_blk00000375 : XORCY
    port map (
      CI => blk00000003_sig000005b5,
      LI => blk00000003_sig000005b6,
      O => blk00000003_sig000005b7
    );
  blk00000003_blk00000374 : XORCY
    port map (
      CI => blk00000003_sig000005b2,
      LI => blk00000003_sig000005b3,
      O => blk00000003_sig000005b4
    );
  blk00000003_blk00000373 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005ad,
      Q => blk00000003_sig000005b1
    );
  blk00000003_blk00000372 : MUXCY
    port map (
      CI => blk00000003_sig000005ae,
      DI => blk00000003_sig00000076,
      S => blk00000003_sig000005af,
      O => blk00000003_sig000005a2
    );
  blk00000003_blk00000371 : XORCY
    port map (
      CI => blk00000003_sig000005ae,
      LI => blk00000003_sig000005af,
      O => blk00000003_sig000005b0
    );
  blk00000003_blk00000370 : MUXCY
    port map (
      CI => blk00000003_sig0000058d,
      DI => blk00000003_sig000005ac,
      S => blk00000003_sig0000058e,
      O => blk00000003_sig000005ad
    );
  blk00000003_blk0000036f : MUXCY
    port map (
      CI => blk00000003_sig000005a2,
      DI => blk00000003_sig000005ab,
      S => blk00000003_sig000005a3,
      O => blk00000003_sig0000059f
    );
  blk00000003_blk0000036e : MUXCY
    port map (
      CI => blk00000003_sig0000059f,
      DI => blk00000003_sig000005aa,
      S => blk00000003_sig000005a0,
      O => blk00000003_sig0000059c
    );
  blk00000003_blk0000036d : MUXCY
    port map (
      CI => blk00000003_sig0000059c,
      DI => blk00000003_sig000005a9,
      S => blk00000003_sig0000059d,
      O => blk00000003_sig00000599
    );
  blk00000003_blk0000036c : MUXCY
    port map (
      CI => blk00000003_sig00000599,
      DI => blk00000003_sig000005a8,
      S => blk00000003_sig0000059a,
      O => blk00000003_sig00000596
    );
  blk00000003_blk0000036b : MUXCY
    port map (
      CI => blk00000003_sig00000596,
      DI => blk00000003_sig000005a7,
      S => blk00000003_sig00000597,
      O => blk00000003_sig00000593
    );
  blk00000003_blk0000036a : MUXCY
    port map (
      CI => blk00000003_sig00000593,
      DI => blk00000003_sig000005a6,
      S => blk00000003_sig00000594,
      O => blk00000003_sig00000590
    );
  blk00000003_blk00000369 : MUXCY
    port map (
      CI => blk00000003_sig00000590,
      DI => blk00000003_sig000005a5,
      S => blk00000003_sig00000591,
      O => blk00000003_sig0000058d
    );
  blk00000003_blk00000368 : XORCY
    port map (
      CI => blk00000003_sig000005a2,
      LI => blk00000003_sig000005a3,
      O => blk00000003_sig000005a4
    );
  blk00000003_blk00000367 : XORCY
    port map (
      CI => blk00000003_sig0000059f,
      LI => blk00000003_sig000005a0,
      O => blk00000003_sig000005a1
    );
  blk00000003_blk00000366 : XORCY
    port map (
      CI => blk00000003_sig0000059c,
      LI => blk00000003_sig0000059d,
      O => blk00000003_sig0000059e
    );
  blk00000003_blk00000365 : XORCY
    port map (
      CI => blk00000003_sig00000599,
      LI => blk00000003_sig0000059a,
      O => blk00000003_sig0000059b
    );
  blk00000003_blk00000364 : XORCY
    port map (
      CI => blk00000003_sig00000596,
      LI => blk00000003_sig00000597,
      O => blk00000003_sig00000598
    );
  blk00000003_blk00000363 : XORCY
    port map (
      CI => blk00000003_sig00000593,
      LI => blk00000003_sig00000594,
      O => blk00000003_sig00000595
    );
  blk00000003_blk00000362 : XORCY
    port map (
      CI => blk00000003_sig00000590,
      LI => blk00000003_sig00000591,
      O => blk00000003_sig00000592
    );
  blk00000003_blk00000361 : XORCY
    port map (
      CI => blk00000003_sig0000058d,
      LI => blk00000003_sig0000058e,
      O => blk00000003_sig0000058f
    );
  blk00000003_blk00000360 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000587,
      Q => blk00000003_sig0000058c
    );
  blk00000003_blk0000035f : MUXCY
    port map (
      CI => blk00000003_sig00000588,
      DI => blk00000003_sig0000058b,
      S => blk00000003_sig00000589,
      O => blk00000003_sig0000057c
    );
  blk00000003_blk0000035e : XORCY
    port map (
      CI => blk00000003_sig00000588,
      LI => blk00000003_sig00000589,
      O => blk00000003_sig0000058a
    );
  blk00000003_blk0000035d : MUXCY
    port map (
      CI => blk00000003_sig00000567,
      DI => blk00000003_sig00000586,
      S => blk00000003_sig00000568,
      O => blk00000003_sig00000587
    );
  blk00000003_blk0000035c : MUXCY
    port map (
      CI => blk00000003_sig0000057c,
      DI => blk00000003_sig00000585,
      S => blk00000003_sig0000057d,
      O => blk00000003_sig00000579
    );
  blk00000003_blk0000035b : MUXCY
    port map (
      CI => blk00000003_sig00000579,
      DI => blk00000003_sig00000584,
      S => blk00000003_sig0000057a,
      O => blk00000003_sig00000576
    );
  blk00000003_blk0000035a : MUXCY
    port map (
      CI => blk00000003_sig00000576,
      DI => blk00000003_sig00000583,
      S => blk00000003_sig00000577,
      O => blk00000003_sig00000573
    );
  blk00000003_blk00000359 : MUXCY
    port map (
      CI => blk00000003_sig00000573,
      DI => blk00000003_sig00000582,
      S => blk00000003_sig00000574,
      O => blk00000003_sig00000570
    );
  blk00000003_blk00000358 : MUXCY
    port map (
      CI => blk00000003_sig00000570,
      DI => blk00000003_sig00000581,
      S => blk00000003_sig00000571,
      O => blk00000003_sig0000056d
    );
  blk00000003_blk00000357 : MUXCY
    port map (
      CI => blk00000003_sig0000056d,
      DI => blk00000003_sig00000580,
      S => blk00000003_sig0000056e,
      O => blk00000003_sig0000056a
    );
  blk00000003_blk00000356 : MUXCY
    port map (
      CI => blk00000003_sig0000056a,
      DI => blk00000003_sig0000057f,
      S => blk00000003_sig0000056b,
      O => blk00000003_sig00000567
    );
  blk00000003_blk00000355 : XORCY
    port map (
      CI => blk00000003_sig0000057c,
      LI => blk00000003_sig0000057d,
      O => blk00000003_sig0000057e
    );
  blk00000003_blk00000354 : XORCY
    port map (
      CI => blk00000003_sig00000579,
      LI => blk00000003_sig0000057a,
      O => blk00000003_sig0000057b
    );
  blk00000003_blk00000353 : XORCY
    port map (
      CI => blk00000003_sig00000576,
      LI => blk00000003_sig00000577,
      O => blk00000003_sig00000578
    );
  blk00000003_blk00000352 : XORCY
    port map (
      CI => blk00000003_sig00000573,
      LI => blk00000003_sig00000574,
      O => blk00000003_sig00000575
    );
  blk00000003_blk00000351 : XORCY
    port map (
      CI => blk00000003_sig00000570,
      LI => blk00000003_sig00000571,
      O => blk00000003_sig00000572
    );
  blk00000003_blk00000350 : XORCY
    port map (
      CI => blk00000003_sig0000056d,
      LI => blk00000003_sig0000056e,
      O => blk00000003_sig0000056f
    );
  blk00000003_blk0000034f : XORCY
    port map (
      CI => blk00000003_sig0000056a,
      LI => blk00000003_sig0000056b,
      O => blk00000003_sig0000056c
    );
  blk00000003_blk0000034e : XORCY
    port map (
      CI => blk00000003_sig00000567,
      LI => blk00000003_sig00000568,
      O => blk00000003_sig00000569
    );
  blk00000003_blk0000034d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000561,
      Q => blk00000003_sig00000566
    );
  blk00000003_blk0000034c : MUXCY
    port map (
      CI => blk00000003_sig00000562,
      DI => blk00000003_sig00000565,
      S => blk00000003_sig00000563,
      O => blk00000003_sig00000556
    );
  blk00000003_blk0000034b : XORCY
    port map (
      CI => blk00000003_sig00000562,
      LI => blk00000003_sig00000563,
      O => blk00000003_sig00000564
    );
  blk00000003_blk0000034a : MUXCY
    port map (
      CI => blk00000003_sig00000541,
      DI => blk00000003_sig00000560,
      S => blk00000003_sig00000542,
      O => blk00000003_sig00000561
    );
  blk00000003_blk00000349 : MUXCY
    port map (
      CI => blk00000003_sig00000556,
      DI => blk00000003_sig0000055f,
      S => blk00000003_sig00000557,
      O => blk00000003_sig00000553
    );
  blk00000003_blk00000348 : MUXCY
    port map (
      CI => blk00000003_sig00000553,
      DI => blk00000003_sig0000055e,
      S => blk00000003_sig00000554,
      O => blk00000003_sig00000550
    );
  blk00000003_blk00000347 : MUXCY
    port map (
      CI => blk00000003_sig00000550,
      DI => blk00000003_sig0000055d,
      S => blk00000003_sig00000551,
      O => blk00000003_sig0000054d
    );
  blk00000003_blk00000346 : MUXCY
    port map (
      CI => blk00000003_sig0000054d,
      DI => blk00000003_sig0000055c,
      S => blk00000003_sig0000054e,
      O => blk00000003_sig0000054a
    );
  blk00000003_blk00000345 : MUXCY
    port map (
      CI => blk00000003_sig0000054a,
      DI => blk00000003_sig0000055b,
      S => blk00000003_sig0000054b,
      O => blk00000003_sig00000547
    );
  blk00000003_blk00000344 : MUXCY
    port map (
      CI => blk00000003_sig00000547,
      DI => blk00000003_sig0000055a,
      S => blk00000003_sig00000548,
      O => blk00000003_sig00000544
    );
  blk00000003_blk00000343 : MUXCY
    port map (
      CI => blk00000003_sig00000544,
      DI => blk00000003_sig00000559,
      S => blk00000003_sig00000545,
      O => blk00000003_sig00000541
    );
  blk00000003_blk00000342 : XORCY
    port map (
      CI => blk00000003_sig00000556,
      LI => blk00000003_sig00000557,
      O => blk00000003_sig00000558
    );
  blk00000003_blk00000341 : XORCY
    port map (
      CI => blk00000003_sig00000553,
      LI => blk00000003_sig00000554,
      O => blk00000003_sig00000555
    );
  blk00000003_blk00000340 : XORCY
    port map (
      CI => blk00000003_sig00000550,
      LI => blk00000003_sig00000551,
      O => blk00000003_sig00000552
    );
  blk00000003_blk0000033f : XORCY
    port map (
      CI => blk00000003_sig0000054d,
      LI => blk00000003_sig0000054e,
      O => blk00000003_sig0000054f
    );
  blk00000003_blk0000033e : XORCY
    port map (
      CI => blk00000003_sig0000054a,
      LI => blk00000003_sig0000054b,
      O => blk00000003_sig0000054c
    );
  blk00000003_blk0000033d : XORCY
    port map (
      CI => blk00000003_sig00000547,
      LI => blk00000003_sig00000548,
      O => blk00000003_sig00000549
    );
  blk00000003_blk0000033c : XORCY
    port map (
      CI => blk00000003_sig00000544,
      LI => blk00000003_sig00000545,
      O => blk00000003_sig00000546
    );
  blk00000003_blk0000033b : XORCY
    port map (
      CI => blk00000003_sig00000541,
      LI => blk00000003_sig00000542,
      O => blk00000003_sig00000543
    );
  blk00000003_blk0000033a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000053b,
      Q => blk00000003_sig00000540
    );
  blk00000003_blk00000339 : MUXCY
    port map (
      CI => blk00000003_sig0000053c,
      DI => blk00000003_sig0000053f,
      S => blk00000003_sig0000053d,
      O => blk00000003_sig00000530
    );
  blk00000003_blk00000338 : XORCY
    port map (
      CI => blk00000003_sig0000053c,
      LI => blk00000003_sig0000053d,
      O => blk00000003_sig0000053e
    );
  blk00000003_blk00000337 : MUXCY
    port map (
      CI => blk00000003_sig0000051b,
      DI => blk00000003_sig0000053a,
      S => blk00000003_sig0000051c,
      O => blk00000003_sig0000053b
    );
  blk00000003_blk00000336 : MUXCY
    port map (
      CI => blk00000003_sig00000530,
      DI => blk00000003_sig00000539,
      S => blk00000003_sig00000531,
      O => blk00000003_sig0000052d
    );
  blk00000003_blk00000335 : MUXCY
    port map (
      CI => blk00000003_sig0000052d,
      DI => blk00000003_sig00000538,
      S => blk00000003_sig0000052e,
      O => blk00000003_sig0000052a
    );
  blk00000003_blk00000334 : MUXCY
    port map (
      CI => blk00000003_sig0000052a,
      DI => blk00000003_sig00000537,
      S => blk00000003_sig0000052b,
      O => blk00000003_sig00000527
    );
  blk00000003_blk00000333 : MUXCY
    port map (
      CI => blk00000003_sig00000527,
      DI => blk00000003_sig00000536,
      S => blk00000003_sig00000528,
      O => blk00000003_sig00000524
    );
  blk00000003_blk00000332 : MUXCY
    port map (
      CI => blk00000003_sig00000524,
      DI => blk00000003_sig00000535,
      S => blk00000003_sig00000525,
      O => blk00000003_sig00000521
    );
  blk00000003_blk00000331 : MUXCY
    port map (
      CI => blk00000003_sig00000521,
      DI => blk00000003_sig00000534,
      S => blk00000003_sig00000522,
      O => blk00000003_sig0000051e
    );
  blk00000003_blk00000330 : MUXCY
    port map (
      CI => blk00000003_sig0000051e,
      DI => blk00000003_sig00000533,
      S => blk00000003_sig0000051f,
      O => blk00000003_sig0000051b
    );
  blk00000003_blk0000032f : XORCY
    port map (
      CI => blk00000003_sig00000530,
      LI => blk00000003_sig00000531,
      O => blk00000003_sig00000532
    );
  blk00000003_blk0000032e : XORCY
    port map (
      CI => blk00000003_sig0000052d,
      LI => blk00000003_sig0000052e,
      O => blk00000003_sig0000052f
    );
  blk00000003_blk0000032d : XORCY
    port map (
      CI => blk00000003_sig0000052a,
      LI => blk00000003_sig0000052b,
      O => blk00000003_sig0000052c
    );
  blk00000003_blk0000032c : XORCY
    port map (
      CI => blk00000003_sig00000527,
      LI => blk00000003_sig00000528,
      O => blk00000003_sig00000529
    );
  blk00000003_blk0000032b : XORCY
    port map (
      CI => blk00000003_sig00000524,
      LI => blk00000003_sig00000525,
      O => blk00000003_sig00000526
    );
  blk00000003_blk0000032a : XORCY
    port map (
      CI => blk00000003_sig00000521,
      LI => blk00000003_sig00000522,
      O => blk00000003_sig00000523
    );
  blk00000003_blk00000329 : XORCY
    port map (
      CI => blk00000003_sig0000051e,
      LI => blk00000003_sig0000051f,
      O => blk00000003_sig00000520
    );
  blk00000003_blk00000328 : XORCY
    port map (
      CI => blk00000003_sig0000051b,
      LI => blk00000003_sig0000051c,
      O => blk00000003_sig0000051d
    );
  blk00000003_blk00000327 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000515,
      Q => blk00000003_sig0000051a
    );
  blk00000003_blk00000326 : MUXCY
    port map (
      CI => blk00000003_sig00000516,
      DI => blk00000003_sig00000519,
      S => blk00000003_sig00000517,
      O => blk00000003_sig0000050a
    );
  blk00000003_blk00000325 : XORCY
    port map (
      CI => blk00000003_sig00000516,
      LI => blk00000003_sig00000517,
      O => blk00000003_sig00000518
    );
  blk00000003_blk00000324 : MUXCY
    port map (
      CI => blk00000003_sig000004f5,
      DI => blk00000003_sig00000514,
      S => blk00000003_sig000004f6,
      O => blk00000003_sig00000515
    );
  blk00000003_blk00000323 : MUXCY
    port map (
      CI => blk00000003_sig0000050a,
      DI => blk00000003_sig00000513,
      S => blk00000003_sig0000050b,
      O => blk00000003_sig00000507
    );
  blk00000003_blk00000322 : MUXCY
    port map (
      CI => blk00000003_sig00000507,
      DI => blk00000003_sig00000512,
      S => blk00000003_sig00000508,
      O => blk00000003_sig00000504
    );
  blk00000003_blk00000321 : MUXCY
    port map (
      CI => blk00000003_sig00000504,
      DI => blk00000003_sig00000511,
      S => blk00000003_sig00000505,
      O => blk00000003_sig00000501
    );
  blk00000003_blk00000320 : MUXCY
    port map (
      CI => blk00000003_sig00000501,
      DI => blk00000003_sig00000510,
      S => blk00000003_sig00000502,
      O => blk00000003_sig000004fe
    );
  blk00000003_blk0000031f : MUXCY
    port map (
      CI => blk00000003_sig000004fe,
      DI => blk00000003_sig0000050f,
      S => blk00000003_sig000004ff,
      O => blk00000003_sig000004fb
    );
  blk00000003_blk0000031e : MUXCY
    port map (
      CI => blk00000003_sig000004fb,
      DI => blk00000003_sig0000050e,
      S => blk00000003_sig000004fc,
      O => blk00000003_sig000004f8
    );
  blk00000003_blk0000031d : MUXCY
    port map (
      CI => blk00000003_sig000004f8,
      DI => blk00000003_sig0000050d,
      S => blk00000003_sig000004f9,
      O => blk00000003_sig000004f5
    );
  blk00000003_blk0000031c : XORCY
    port map (
      CI => blk00000003_sig0000050a,
      LI => blk00000003_sig0000050b,
      O => blk00000003_sig0000050c
    );
  blk00000003_blk0000031b : XORCY
    port map (
      CI => blk00000003_sig00000507,
      LI => blk00000003_sig00000508,
      O => blk00000003_sig00000509
    );
  blk00000003_blk0000031a : XORCY
    port map (
      CI => blk00000003_sig00000504,
      LI => blk00000003_sig00000505,
      O => blk00000003_sig00000506
    );
  blk00000003_blk00000319 : XORCY
    port map (
      CI => blk00000003_sig00000501,
      LI => blk00000003_sig00000502,
      O => blk00000003_sig00000503
    );
  blk00000003_blk00000318 : XORCY
    port map (
      CI => blk00000003_sig000004fe,
      LI => blk00000003_sig000004ff,
      O => blk00000003_sig00000500
    );
  blk00000003_blk00000317 : XORCY
    port map (
      CI => blk00000003_sig000004fb,
      LI => blk00000003_sig000004fc,
      O => blk00000003_sig000004fd
    );
  blk00000003_blk00000316 : XORCY
    port map (
      CI => blk00000003_sig000004f8,
      LI => blk00000003_sig000004f9,
      O => blk00000003_sig000004fa
    );
  blk00000003_blk00000315 : XORCY
    port map (
      CI => blk00000003_sig000004f5,
      LI => blk00000003_sig000004f6,
      O => blk00000003_sig000004f7
    );
  blk00000003_blk00000314 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004ef,
      Q => blk00000003_sig000004f4
    );
  blk00000003_blk00000313 : MUXCY
    port map (
      CI => blk00000003_sig000004f0,
      DI => blk00000003_sig000004f3,
      S => blk00000003_sig000004f1,
      O => blk00000003_sig000004e4
    );
  blk00000003_blk00000312 : XORCY
    port map (
      CI => blk00000003_sig000004f0,
      LI => blk00000003_sig000004f1,
      O => blk00000003_sig000004f2
    );
  blk00000003_blk00000311 : MUXCY
    port map (
      CI => blk00000003_sig000004cf,
      DI => blk00000003_sig000004ee,
      S => blk00000003_sig000004d0,
      O => blk00000003_sig000004ef
    );
  blk00000003_blk00000310 : MUXCY
    port map (
      CI => blk00000003_sig000004e4,
      DI => blk00000003_sig000004ed,
      S => blk00000003_sig000004e5,
      O => blk00000003_sig000004e1
    );
  blk00000003_blk0000030f : MUXCY
    port map (
      CI => blk00000003_sig000004e1,
      DI => blk00000003_sig000004ec,
      S => blk00000003_sig000004e2,
      O => blk00000003_sig000004de
    );
  blk00000003_blk0000030e : MUXCY
    port map (
      CI => blk00000003_sig000004de,
      DI => blk00000003_sig000004eb,
      S => blk00000003_sig000004df,
      O => blk00000003_sig000004db
    );
  blk00000003_blk0000030d : MUXCY
    port map (
      CI => blk00000003_sig000004db,
      DI => blk00000003_sig000004ea,
      S => blk00000003_sig000004dc,
      O => blk00000003_sig000004d8
    );
  blk00000003_blk0000030c : MUXCY
    port map (
      CI => blk00000003_sig000004d8,
      DI => blk00000003_sig000004e9,
      S => blk00000003_sig000004d9,
      O => blk00000003_sig000004d5
    );
  blk00000003_blk0000030b : MUXCY
    port map (
      CI => blk00000003_sig000004d5,
      DI => blk00000003_sig000004e8,
      S => blk00000003_sig000004d6,
      O => blk00000003_sig000004d2
    );
  blk00000003_blk0000030a : MUXCY
    port map (
      CI => blk00000003_sig000004d2,
      DI => blk00000003_sig000004e7,
      S => blk00000003_sig000004d3,
      O => blk00000003_sig000004cf
    );
  blk00000003_blk00000309 : XORCY
    port map (
      CI => blk00000003_sig000004e4,
      LI => blk00000003_sig000004e5,
      O => blk00000003_sig000004e6
    );
  blk00000003_blk00000308 : XORCY
    port map (
      CI => blk00000003_sig000004e1,
      LI => blk00000003_sig000004e2,
      O => blk00000003_sig000004e3
    );
  blk00000003_blk00000307 : XORCY
    port map (
      CI => blk00000003_sig000004de,
      LI => blk00000003_sig000004df,
      O => blk00000003_sig000004e0
    );
  blk00000003_blk00000306 : XORCY
    port map (
      CI => blk00000003_sig000004db,
      LI => blk00000003_sig000004dc,
      O => blk00000003_sig000004dd
    );
  blk00000003_blk00000305 : XORCY
    port map (
      CI => blk00000003_sig000004d8,
      LI => blk00000003_sig000004d9,
      O => blk00000003_sig000004da
    );
  blk00000003_blk00000304 : XORCY
    port map (
      CI => blk00000003_sig000004d5,
      LI => blk00000003_sig000004d6,
      O => blk00000003_sig000004d7
    );
  blk00000003_blk00000303 : XORCY
    port map (
      CI => blk00000003_sig000004d2,
      LI => blk00000003_sig000004d3,
      O => blk00000003_sig000004d4
    );
  blk00000003_blk00000302 : XORCY
    port map (
      CI => blk00000003_sig000004cf,
      LI => blk00000003_sig000004d0,
      O => blk00000003_sig000004d1
    );
  blk00000003_blk00000301 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004c9,
      Q => blk00000003_sig000004ce
    );
  blk00000003_blk00000300 : MUXCY
    port map (
      CI => blk00000003_sig000004ca,
      DI => blk00000003_sig000004cd,
      S => blk00000003_sig000004cb,
      O => blk00000003_sig000004be
    );
  blk00000003_blk000002ff : XORCY
    port map (
      CI => blk00000003_sig000004ca,
      LI => blk00000003_sig000004cb,
      O => blk00000003_sig000004cc
    );
  blk00000003_blk000002fe : MUXCY
    port map (
      CI => blk00000003_sig000004a9,
      DI => blk00000003_sig000004c8,
      S => blk00000003_sig000004aa,
      O => blk00000003_sig000004c9
    );
  blk00000003_blk000002fd : MUXCY
    port map (
      CI => blk00000003_sig000004be,
      DI => blk00000003_sig000004c7,
      S => blk00000003_sig000004bf,
      O => blk00000003_sig000004bb
    );
  blk00000003_blk000002fc : MUXCY
    port map (
      CI => blk00000003_sig000004bb,
      DI => blk00000003_sig000004c6,
      S => blk00000003_sig000004bc,
      O => blk00000003_sig000004b8
    );
  blk00000003_blk000002fb : MUXCY
    port map (
      CI => blk00000003_sig000004b8,
      DI => blk00000003_sig000004c5,
      S => blk00000003_sig000004b9,
      O => blk00000003_sig000004b5
    );
  blk00000003_blk000002fa : MUXCY
    port map (
      CI => blk00000003_sig000004b5,
      DI => blk00000003_sig000004c4,
      S => blk00000003_sig000004b6,
      O => blk00000003_sig000004b2
    );
  blk00000003_blk000002f9 : MUXCY
    port map (
      CI => blk00000003_sig000004b2,
      DI => blk00000003_sig000004c3,
      S => blk00000003_sig000004b3,
      O => blk00000003_sig000004af
    );
  blk00000003_blk000002f8 : MUXCY
    port map (
      CI => blk00000003_sig000004af,
      DI => blk00000003_sig000004c2,
      S => blk00000003_sig000004b0,
      O => blk00000003_sig000004ac
    );
  blk00000003_blk000002f7 : MUXCY
    port map (
      CI => blk00000003_sig000004ac,
      DI => blk00000003_sig000004c1,
      S => blk00000003_sig000004ad,
      O => blk00000003_sig000004a9
    );
  blk00000003_blk000002f6 : XORCY
    port map (
      CI => blk00000003_sig000004be,
      LI => blk00000003_sig000004bf,
      O => blk00000003_sig000004c0
    );
  blk00000003_blk000002f5 : XORCY
    port map (
      CI => blk00000003_sig000004bb,
      LI => blk00000003_sig000004bc,
      O => blk00000003_sig000004bd
    );
  blk00000003_blk000002f4 : XORCY
    port map (
      CI => blk00000003_sig000004b8,
      LI => blk00000003_sig000004b9,
      O => blk00000003_sig000004ba
    );
  blk00000003_blk000002f3 : XORCY
    port map (
      CI => blk00000003_sig000004b5,
      LI => blk00000003_sig000004b6,
      O => blk00000003_sig000004b7
    );
  blk00000003_blk000002f2 : XORCY
    port map (
      CI => blk00000003_sig000004b2,
      LI => blk00000003_sig000004b3,
      O => blk00000003_sig000004b4
    );
  blk00000003_blk000002f1 : XORCY
    port map (
      CI => blk00000003_sig000004af,
      LI => blk00000003_sig000004b0,
      O => blk00000003_sig000004b1
    );
  blk00000003_blk000002f0 : XORCY
    port map (
      CI => blk00000003_sig000004ac,
      LI => blk00000003_sig000004ad,
      O => blk00000003_sig000004ae
    );
  blk00000003_blk000002ef : XORCY
    port map (
      CI => blk00000003_sig000004a9,
      LI => blk00000003_sig000004aa,
      O => blk00000003_sig000004ab
    );
  blk00000003_blk000002ee : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004a3,
      Q => blk00000003_sig000004a8
    );
  blk00000003_blk000002ed : MUXCY
    port map (
      CI => blk00000003_sig000004a4,
      DI => blk00000003_sig000004a7,
      S => blk00000003_sig000004a5,
      O => blk00000003_sig00000498
    );
  blk00000003_blk000002ec : XORCY
    port map (
      CI => blk00000003_sig000004a4,
      LI => blk00000003_sig000004a5,
      O => blk00000003_sig000004a6
    );
  blk00000003_blk000002eb : MUXCY
    port map (
      CI => blk00000003_sig00000483,
      DI => blk00000003_sig000004a2,
      S => blk00000003_sig00000484,
      O => blk00000003_sig000004a3
    );
  blk00000003_blk000002ea : MUXCY
    port map (
      CI => blk00000003_sig00000498,
      DI => blk00000003_sig000004a1,
      S => blk00000003_sig00000499,
      O => blk00000003_sig00000495
    );
  blk00000003_blk000002e9 : MUXCY
    port map (
      CI => blk00000003_sig00000495,
      DI => blk00000003_sig000004a0,
      S => blk00000003_sig00000496,
      O => blk00000003_sig00000492
    );
  blk00000003_blk000002e8 : MUXCY
    port map (
      CI => blk00000003_sig00000492,
      DI => blk00000003_sig0000049f,
      S => blk00000003_sig00000493,
      O => blk00000003_sig0000048f
    );
  blk00000003_blk000002e7 : MUXCY
    port map (
      CI => blk00000003_sig0000048f,
      DI => blk00000003_sig0000049e,
      S => blk00000003_sig00000490,
      O => blk00000003_sig0000048c
    );
  blk00000003_blk000002e6 : MUXCY
    port map (
      CI => blk00000003_sig0000048c,
      DI => blk00000003_sig0000049d,
      S => blk00000003_sig0000048d,
      O => blk00000003_sig00000489
    );
  blk00000003_blk000002e5 : MUXCY
    port map (
      CI => blk00000003_sig00000489,
      DI => blk00000003_sig0000049c,
      S => blk00000003_sig0000048a,
      O => blk00000003_sig00000486
    );
  blk00000003_blk000002e4 : MUXCY
    port map (
      CI => blk00000003_sig00000486,
      DI => blk00000003_sig0000049b,
      S => blk00000003_sig00000487,
      O => blk00000003_sig00000483
    );
  blk00000003_blk000002e3 : XORCY
    port map (
      CI => blk00000003_sig00000498,
      LI => blk00000003_sig00000499,
      O => blk00000003_sig0000049a
    );
  blk00000003_blk000002e2 : XORCY
    port map (
      CI => blk00000003_sig00000495,
      LI => blk00000003_sig00000496,
      O => blk00000003_sig00000497
    );
  blk00000003_blk000002e1 : XORCY
    port map (
      CI => blk00000003_sig00000492,
      LI => blk00000003_sig00000493,
      O => blk00000003_sig00000494
    );
  blk00000003_blk000002e0 : XORCY
    port map (
      CI => blk00000003_sig0000048f,
      LI => blk00000003_sig00000490,
      O => blk00000003_sig00000491
    );
  blk00000003_blk000002df : XORCY
    port map (
      CI => blk00000003_sig0000048c,
      LI => blk00000003_sig0000048d,
      O => blk00000003_sig0000048e
    );
  blk00000003_blk000002de : XORCY
    port map (
      CI => blk00000003_sig00000489,
      LI => blk00000003_sig0000048a,
      O => blk00000003_sig0000048b
    );
  blk00000003_blk000002dd : XORCY
    port map (
      CI => blk00000003_sig00000486,
      LI => blk00000003_sig00000487,
      O => blk00000003_sig00000488
    );
  blk00000003_blk000002dc : XORCY
    port map (
      CI => blk00000003_sig00000483,
      LI => blk00000003_sig00000484,
      O => blk00000003_sig00000485
    );
  blk00000003_blk000002db : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000047d,
      Q => blk00000003_sig00000482
    );
  blk00000003_blk000002da : MUXCY
    port map (
      CI => blk00000003_sig0000047e,
      DI => blk00000003_sig00000481,
      S => blk00000003_sig0000047f,
      O => blk00000003_sig00000472
    );
  blk00000003_blk000002d9 : XORCY
    port map (
      CI => blk00000003_sig0000047e,
      LI => blk00000003_sig0000047f,
      O => blk00000003_sig00000480
    );
  blk00000003_blk000002d8 : MUXCY
    port map (
      CI => blk00000003_sig0000045d,
      DI => blk00000003_sig0000047c,
      S => blk00000003_sig0000045e,
      O => blk00000003_sig0000047d
    );
  blk00000003_blk000002d7 : MUXCY
    port map (
      CI => blk00000003_sig00000472,
      DI => blk00000003_sig0000047b,
      S => blk00000003_sig00000473,
      O => blk00000003_sig0000046f
    );
  blk00000003_blk000002d6 : MUXCY
    port map (
      CI => blk00000003_sig0000046f,
      DI => blk00000003_sig0000047a,
      S => blk00000003_sig00000470,
      O => blk00000003_sig0000046c
    );
  blk00000003_blk000002d5 : MUXCY
    port map (
      CI => blk00000003_sig0000046c,
      DI => blk00000003_sig00000479,
      S => blk00000003_sig0000046d,
      O => blk00000003_sig00000469
    );
  blk00000003_blk000002d4 : MUXCY
    port map (
      CI => blk00000003_sig00000469,
      DI => blk00000003_sig00000478,
      S => blk00000003_sig0000046a,
      O => blk00000003_sig00000466
    );
  blk00000003_blk000002d3 : MUXCY
    port map (
      CI => blk00000003_sig00000466,
      DI => blk00000003_sig00000477,
      S => blk00000003_sig00000467,
      O => blk00000003_sig00000463
    );
  blk00000003_blk000002d2 : MUXCY
    port map (
      CI => blk00000003_sig00000463,
      DI => blk00000003_sig00000476,
      S => blk00000003_sig00000464,
      O => blk00000003_sig00000460
    );
  blk00000003_blk000002d1 : MUXCY
    port map (
      CI => blk00000003_sig00000460,
      DI => blk00000003_sig00000475,
      S => blk00000003_sig00000461,
      O => blk00000003_sig0000045d
    );
  blk00000003_blk000002d0 : XORCY
    port map (
      CI => blk00000003_sig00000472,
      LI => blk00000003_sig00000473,
      O => blk00000003_sig00000474
    );
  blk00000003_blk000002cf : XORCY
    port map (
      CI => blk00000003_sig0000046f,
      LI => blk00000003_sig00000470,
      O => blk00000003_sig00000471
    );
  blk00000003_blk000002ce : XORCY
    port map (
      CI => blk00000003_sig0000046c,
      LI => blk00000003_sig0000046d,
      O => blk00000003_sig0000046e
    );
  blk00000003_blk000002cd : XORCY
    port map (
      CI => blk00000003_sig00000469,
      LI => blk00000003_sig0000046a,
      O => blk00000003_sig0000046b
    );
  blk00000003_blk000002cc : XORCY
    port map (
      CI => blk00000003_sig00000466,
      LI => blk00000003_sig00000467,
      O => blk00000003_sig00000468
    );
  blk00000003_blk000002cb : XORCY
    port map (
      CI => blk00000003_sig00000463,
      LI => blk00000003_sig00000464,
      O => blk00000003_sig00000465
    );
  blk00000003_blk000002ca : XORCY
    port map (
      CI => blk00000003_sig00000460,
      LI => blk00000003_sig00000461,
      O => blk00000003_sig00000462
    );
  blk00000003_blk000002c9 : XORCY
    port map (
      CI => blk00000003_sig0000045d,
      LI => blk00000003_sig0000045e,
      O => blk00000003_sig0000045f
    );
  blk00000003_blk000002c8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000457,
      Q => blk00000003_sig0000045c
    );
  blk00000003_blk000002c7 : MUXCY
    port map (
      CI => blk00000003_sig00000458,
      DI => blk00000003_sig0000045b,
      S => blk00000003_sig00000459,
      O => blk00000003_sig0000044c
    );
  blk00000003_blk000002c6 : XORCY
    port map (
      CI => blk00000003_sig00000458,
      LI => blk00000003_sig00000459,
      O => blk00000003_sig0000045a
    );
  blk00000003_blk000002c5 : MUXCY
    port map (
      CI => blk00000003_sig00000437,
      DI => blk00000003_sig00000456,
      S => blk00000003_sig00000438,
      O => blk00000003_sig00000457
    );
  blk00000003_blk000002c4 : MUXCY
    port map (
      CI => blk00000003_sig0000044c,
      DI => blk00000003_sig00000455,
      S => blk00000003_sig0000044d,
      O => blk00000003_sig00000449
    );
  blk00000003_blk000002c3 : MUXCY
    port map (
      CI => blk00000003_sig00000449,
      DI => blk00000003_sig00000454,
      S => blk00000003_sig0000044a,
      O => blk00000003_sig00000446
    );
  blk00000003_blk000002c2 : MUXCY
    port map (
      CI => blk00000003_sig00000446,
      DI => blk00000003_sig00000453,
      S => blk00000003_sig00000447,
      O => blk00000003_sig00000443
    );
  blk00000003_blk000002c1 : MUXCY
    port map (
      CI => blk00000003_sig00000443,
      DI => blk00000003_sig00000452,
      S => blk00000003_sig00000444,
      O => blk00000003_sig00000440
    );
  blk00000003_blk000002c0 : MUXCY
    port map (
      CI => blk00000003_sig00000440,
      DI => blk00000003_sig00000451,
      S => blk00000003_sig00000441,
      O => blk00000003_sig0000043d
    );
  blk00000003_blk000002bf : MUXCY
    port map (
      CI => blk00000003_sig0000043d,
      DI => blk00000003_sig00000450,
      S => blk00000003_sig0000043e,
      O => blk00000003_sig0000043a
    );
  blk00000003_blk000002be : MUXCY
    port map (
      CI => blk00000003_sig0000043a,
      DI => blk00000003_sig0000044f,
      S => blk00000003_sig0000043b,
      O => blk00000003_sig00000437
    );
  blk00000003_blk000002bd : XORCY
    port map (
      CI => blk00000003_sig0000044c,
      LI => blk00000003_sig0000044d,
      O => blk00000003_sig0000044e
    );
  blk00000003_blk000002bc : XORCY
    port map (
      CI => blk00000003_sig00000449,
      LI => blk00000003_sig0000044a,
      O => blk00000003_sig0000044b
    );
  blk00000003_blk000002bb : XORCY
    port map (
      CI => blk00000003_sig00000446,
      LI => blk00000003_sig00000447,
      O => blk00000003_sig00000448
    );
  blk00000003_blk000002ba : XORCY
    port map (
      CI => blk00000003_sig00000443,
      LI => blk00000003_sig00000444,
      O => blk00000003_sig00000445
    );
  blk00000003_blk000002b9 : XORCY
    port map (
      CI => blk00000003_sig00000440,
      LI => blk00000003_sig00000441,
      O => blk00000003_sig00000442
    );
  blk00000003_blk000002b8 : XORCY
    port map (
      CI => blk00000003_sig0000043d,
      LI => blk00000003_sig0000043e,
      O => blk00000003_sig0000043f
    );
  blk00000003_blk000002b7 : XORCY
    port map (
      CI => blk00000003_sig0000043a,
      LI => blk00000003_sig0000043b,
      O => blk00000003_sig0000043c
    );
  blk00000003_blk000002b6 : XORCY
    port map (
      CI => blk00000003_sig00000437,
      LI => blk00000003_sig00000438,
      O => blk00000003_sig00000439
    );
  blk00000003_blk000002b5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000431,
      Q => blk00000003_sig00000436
    );
  blk00000003_blk000002b4 : MUXCY
    port map (
      CI => blk00000003_sig00000432,
      DI => blk00000003_sig00000435,
      S => blk00000003_sig00000433,
      O => blk00000003_sig00000426
    );
  blk00000003_blk000002b3 : XORCY
    port map (
      CI => blk00000003_sig00000432,
      LI => blk00000003_sig00000433,
      O => blk00000003_sig00000434
    );
  blk00000003_blk000002b2 : MUXCY
    port map (
      CI => blk00000003_sig00000411,
      DI => blk00000003_sig00000430,
      S => blk00000003_sig00000412,
      O => blk00000003_sig00000431
    );
  blk00000003_blk000002b1 : MUXCY
    port map (
      CI => blk00000003_sig00000426,
      DI => blk00000003_sig0000042f,
      S => blk00000003_sig00000427,
      O => blk00000003_sig00000423
    );
  blk00000003_blk000002b0 : MUXCY
    port map (
      CI => blk00000003_sig00000423,
      DI => blk00000003_sig0000042e,
      S => blk00000003_sig00000424,
      O => blk00000003_sig00000420
    );
  blk00000003_blk000002af : MUXCY
    port map (
      CI => blk00000003_sig00000420,
      DI => blk00000003_sig0000042d,
      S => blk00000003_sig00000421,
      O => blk00000003_sig0000041d
    );
  blk00000003_blk000002ae : MUXCY
    port map (
      CI => blk00000003_sig0000041d,
      DI => blk00000003_sig0000042c,
      S => blk00000003_sig0000041e,
      O => blk00000003_sig0000041a
    );
  blk00000003_blk000002ad : MUXCY
    port map (
      CI => blk00000003_sig0000041a,
      DI => blk00000003_sig0000042b,
      S => blk00000003_sig0000041b,
      O => blk00000003_sig00000417
    );
  blk00000003_blk000002ac : MUXCY
    port map (
      CI => blk00000003_sig00000417,
      DI => blk00000003_sig0000042a,
      S => blk00000003_sig00000418,
      O => blk00000003_sig00000414
    );
  blk00000003_blk000002ab : MUXCY
    port map (
      CI => blk00000003_sig00000414,
      DI => blk00000003_sig00000429,
      S => blk00000003_sig00000415,
      O => blk00000003_sig00000411
    );
  blk00000003_blk000002aa : XORCY
    port map (
      CI => blk00000003_sig00000426,
      LI => blk00000003_sig00000427,
      O => blk00000003_sig00000428
    );
  blk00000003_blk000002a9 : XORCY
    port map (
      CI => blk00000003_sig00000423,
      LI => blk00000003_sig00000424,
      O => blk00000003_sig00000425
    );
  blk00000003_blk000002a8 : XORCY
    port map (
      CI => blk00000003_sig00000420,
      LI => blk00000003_sig00000421,
      O => blk00000003_sig00000422
    );
  blk00000003_blk000002a7 : XORCY
    port map (
      CI => blk00000003_sig0000041d,
      LI => blk00000003_sig0000041e,
      O => blk00000003_sig0000041f
    );
  blk00000003_blk000002a6 : XORCY
    port map (
      CI => blk00000003_sig0000041a,
      LI => blk00000003_sig0000041b,
      O => blk00000003_sig0000041c
    );
  blk00000003_blk000002a5 : XORCY
    port map (
      CI => blk00000003_sig00000417,
      LI => blk00000003_sig00000418,
      O => blk00000003_sig00000419
    );
  blk00000003_blk000002a4 : XORCY
    port map (
      CI => blk00000003_sig00000414,
      LI => blk00000003_sig00000415,
      O => blk00000003_sig00000416
    );
  blk00000003_blk000002a3 : XORCY
    port map (
      CI => blk00000003_sig00000411,
      LI => blk00000003_sig00000412,
      O => blk00000003_sig00000413
    );
  blk00000003_blk000002a2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000040b,
      Q => blk00000003_sig00000410
    );
  blk00000003_blk000002a1 : MUXCY
    port map (
      CI => blk00000003_sig0000040c,
      DI => blk00000003_sig0000040f,
      S => blk00000003_sig0000040d,
      O => blk00000003_sig00000400
    );
  blk00000003_blk000002a0 : XORCY
    port map (
      CI => blk00000003_sig0000040c,
      LI => blk00000003_sig0000040d,
      O => blk00000003_sig0000040e
    );
  blk00000003_blk0000029f : MUXCY
    port map (
      CI => blk00000003_sig000003eb,
      DI => blk00000003_sig0000040a,
      S => blk00000003_sig000003ec,
      O => blk00000003_sig0000040b
    );
  blk00000003_blk0000029e : MUXCY
    port map (
      CI => blk00000003_sig00000400,
      DI => blk00000003_sig00000409,
      S => blk00000003_sig00000401,
      O => blk00000003_sig000003fd
    );
  blk00000003_blk0000029d : MUXCY
    port map (
      CI => blk00000003_sig000003fd,
      DI => blk00000003_sig00000408,
      S => blk00000003_sig000003fe,
      O => blk00000003_sig000003fa
    );
  blk00000003_blk0000029c : MUXCY
    port map (
      CI => blk00000003_sig000003fa,
      DI => blk00000003_sig00000407,
      S => blk00000003_sig000003fb,
      O => blk00000003_sig000003f7
    );
  blk00000003_blk0000029b : MUXCY
    port map (
      CI => blk00000003_sig000003f7,
      DI => blk00000003_sig00000406,
      S => blk00000003_sig000003f8,
      O => blk00000003_sig000003f4
    );
  blk00000003_blk0000029a : MUXCY
    port map (
      CI => blk00000003_sig000003f4,
      DI => blk00000003_sig00000405,
      S => blk00000003_sig000003f5,
      O => blk00000003_sig000003f1
    );
  blk00000003_blk00000299 : MUXCY
    port map (
      CI => blk00000003_sig000003f1,
      DI => blk00000003_sig00000404,
      S => blk00000003_sig000003f2,
      O => blk00000003_sig000003ee
    );
  blk00000003_blk00000298 : MUXCY
    port map (
      CI => blk00000003_sig000003ee,
      DI => blk00000003_sig00000403,
      S => blk00000003_sig000003ef,
      O => blk00000003_sig000003eb
    );
  blk00000003_blk00000297 : XORCY
    port map (
      CI => blk00000003_sig00000400,
      LI => blk00000003_sig00000401,
      O => blk00000003_sig00000402
    );
  blk00000003_blk00000296 : XORCY
    port map (
      CI => blk00000003_sig000003fd,
      LI => blk00000003_sig000003fe,
      O => blk00000003_sig000003ff
    );
  blk00000003_blk00000295 : XORCY
    port map (
      CI => blk00000003_sig000003fa,
      LI => blk00000003_sig000003fb,
      O => blk00000003_sig000003fc
    );
  blk00000003_blk00000294 : XORCY
    port map (
      CI => blk00000003_sig000003f7,
      LI => blk00000003_sig000003f8,
      O => blk00000003_sig000003f9
    );
  blk00000003_blk00000293 : XORCY
    port map (
      CI => blk00000003_sig000003f4,
      LI => blk00000003_sig000003f5,
      O => blk00000003_sig000003f6
    );
  blk00000003_blk00000292 : XORCY
    port map (
      CI => blk00000003_sig000003f1,
      LI => blk00000003_sig000003f2,
      O => blk00000003_sig000003f3
    );
  blk00000003_blk00000291 : XORCY
    port map (
      CI => blk00000003_sig000003ee,
      LI => blk00000003_sig000003ef,
      O => blk00000003_sig000003f0
    );
  blk00000003_blk00000290 : XORCY
    port map (
      CI => blk00000003_sig000003eb,
      LI => blk00000003_sig000003ec,
      O => blk00000003_sig000003ed
    );
  blk00000003_blk0000028f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003e5,
      Q => blk00000003_sig000003ea
    );
  blk00000003_blk0000028e : MUXCY
    port map (
      CI => blk00000003_sig000003e6,
      DI => blk00000003_sig000003e9,
      S => blk00000003_sig000003e7,
      O => blk00000003_sig000003da
    );
  blk00000003_blk0000028d : XORCY
    port map (
      CI => blk00000003_sig000003e6,
      LI => blk00000003_sig000003e7,
      O => blk00000003_sig000003e8
    );
  blk00000003_blk0000028c : MUXCY
    port map (
      CI => blk00000003_sig000003c5,
      DI => blk00000003_sig000003e4,
      S => blk00000003_sig000003c6,
      O => blk00000003_sig000003e5
    );
  blk00000003_blk0000028b : MUXCY
    port map (
      CI => blk00000003_sig000003da,
      DI => blk00000003_sig000003e3,
      S => blk00000003_sig000003db,
      O => blk00000003_sig000003d7
    );
  blk00000003_blk0000028a : MUXCY
    port map (
      CI => blk00000003_sig000003d7,
      DI => blk00000003_sig000003e2,
      S => blk00000003_sig000003d8,
      O => blk00000003_sig000003d4
    );
  blk00000003_blk00000289 : MUXCY
    port map (
      CI => blk00000003_sig000003d4,
      DI => blk00000003_sig000003e1,
      S => blk00000003_sig000003d5,
      O => blk00000003_sig000003d1
    );
  blk00000003_blk00000288 : MUXCY
    port map (
      CI => blk00000003_sig000003d1,
      DI => blk00000003_sig000003e0,
      S => blk00000003_sig000003d2,
      O => blk00000003_sig000003ce
    );
  blk00000003_blk00000287 : MUXCY
    port map (
      CI => blk00000003_sig000003ce,
      DI => blk00000003_sig000003df,
      S => blk00000003_sig000003cf,
      O => blk00000003_sig000003cb
    );
  blk00000003_blk00000286 : MUXCY
    port map (
      CI => blk00000003_sig000003cb,
      DI => blk00000003_sig000003de,
      S => blk00000003_sig000003cc,
      O => blk00000003_sig000003c8
    );
  blk00000003_blk00000285 : MUXCY
    port map (
      CI => blk00000003_sig000003c8,
      DI => blk00000003_sig000003dd,
      S => blk00000003_sig000003c9,
      O => blk00000003_sig000003c5
    );
  blk00000003_blk00000284 : XORCY
    port map (
      CI => blk00000003_sig000003da,
      LI => blk00000003_sig000003db,
      O => blk00000003_sig000003dc
    );
  blk00000003_blk00000283 : XORCY
    port map (
      CI => blk00000003_sig000003d7,
      LI => blk00000003_sig000003d8,
      O => blk00000003_sig000003d9
    );
  blk00000003_blk00000282 : XORCY
    port map (
      CI => blk00000003_sig000003d4,
      LI => blk00000003_sig000003d5,
      O => blk00000003_sig000003d6
    );
  blk00000003_blk00000281 : XORCY
    port map (
      CI => blk00000003_sig000003d1,
      LI => blk00000003_sig000003d2,
      O => blk00000003_sig000003d3
    );
  blk00000003_blk00000280 : XORCY
    port map (
      CI => blk00000003_sig000003ce,
      LI => blk00000003_sig000003cf,
      O => blk00000003_sig000003d0
    );
  blk00000003_blk0000027f : XORCY
    port map (
      CI => blk00000003_sig000003cb,
      LI => blk00000003_sig000003cc,
      O => blk00000003_sig000003cd
    );
  blk00000003_blk0000027e : XORCY
    port map (
      CI => blk00000003_sig000003c8,
      LI => blk00000003_sig000003c9,
      O => blk00000003_sig000003ca
    );
  blk00000003_blk0000027d : XORCY
    port map (
      CI => blk00000003_sig000003c5,
      LI => blk00000003_sig000003c6,
      O => blk00000003_sig000003c7
    );
  blk00000003_blk0000027c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003bf,
      Q => blk00000003_sig000003c4
    );
  blk00000003_blk0000027b : MUXCY
    port map (
      CI => blk00000003_sig000003c0,
      DI => blk00000003_sig000003c3,
      S => blk00000003_sig000003c1,
      O => blk00000003_sig000003b4
    );
  blk00000003_blk0000027a : XORCY
    port map (
      CI => blk00000003_sig000003c0,
      LI => blk00000003_sig000003c1,
      O => blk00000003_sig000003c2
    );
  blk00000003_blk00000279 : MUXCY
    port map (
      CI => blk00000003_sig0000039f,
      DI => blk00000003_sig000003be,
      S => blk00000003_sig000003a0,
      O => blk00000003_sig000003bf
    );
  blk00000003_blk00000278 : MUXCY
    port map (
      CI => blk00000003_sig000003b4,
      DI => blk00000003_sig000003bd,
      S => blk00000003_sig000003b5,
      O => blk00000003_sig000003b1
    );
  blk00000003_blk00000277 : MUXCY
    port map (
      CI => blk00000003_sig000003b1,
      DI => blk00000003_sig000003bc,
      S => blk00000003_sig000003b2,
      O => blk00000003_sig000003ae
    );
  blk00000003_blk00000276 : MUXCY
    port map (
      CI => blk00000003_sig000003ae,
      DI => blk00000003_sig000003bb,
      S => blk00000003_sig000003af,
      O => blk00000003_sig000003ab
    );
  blk00000003_blk00000275 : MUXCY
    port map (
      CI => blk00000003_sig000003ab,
      DI => blk00000003_sig000003ba,
      S => blk00000003_sig000003ac,
      O => blk00000003_sig000003a8
    );
  blk00000003_blk00000274 : MUXCY
    port map (
      CI => blk00000003_sig000003a8,
      DI => blk00000003_sig000003b9,
      S => blk00000003_sig000003a9,
      O => blk00000003_sig000003a5
    );
  blk00000003_blk00000273 : MUXCY
    port map (
      CI => blk00000003_sig000003a5,
      DI => blk00000003_sig000003b8,
      S => blk00000003_sig000003a6,
      O => blk00000003_sig000003a2
    );
  blk00000003_blk00000272 : MUXCY
    port map (
      CI => blk00000003_sig000003a2,
      DI => blk00000003_sig000003b7,
      S => blk00000003_sig000003a3,
      O => blk00000003_sig0000039f
    );
  blk00000003_blk00000271 : XORCY
    port map (
      CI => blk00000003_sig000003b4,
      LI => blk00000003_sig000003b5,
      O => blk00000003_sig000003b6
    );
  blk00000003_blk00000270 : XORCY
    port map (
      CI => blk00000003_sig000003b1,
      LI => blk00000003_sig000003b2,
      O => blk00000003_sig000003b3
    );
  blk00000003_blk0000026f : XORCY
    port map (
      CI => blk00000003_sig000003ae,
      LI => blk00000003_sig000003af,
      O => blk00000003_sig000003b0
    );
  blk00000003_blk0000026e : XORCY
    port map (
      CI => blk00000003_sig000003ab,
      LI => blk00000003_sig000003ac,
      O => blk00000003_sig000003ad
    );
  blk00000003_blk0000026d : XORCY
    port map (
      CI => blk00000003_sig000003a8,
      LI => blk00000003_sig000003a9,
      O => blk00000003_sig000003aa
    );
  blk00000003_blk0000026c : XORCY
    port map (
      CI => blk00000003_sig000003a5,
      LI => blk00000003_sig000003a6,
      O => blk00000003_sig000003a7
    );
  blk00000003_blk0000026b : XORCY
    port map (
      CI => blk00000003_sig000003a2,
      LI => blk00000003_sig000003a3,
      O => blk00000003_sig000003a4
    );
  blk00000003_blk0000026a : XORCY
    port map (
      CI => blk00000003_sig0000039f,
      LI => blk00000003_sig000003a0,
      O => blk00000003_sig000003a1
    );
  blk00000003_blk00000269 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000399,
      Q => blk00000003_sig0000039e
    );
  blk00000003_blk00000268 : MUXCY
    port map (
      CI => blk00000003_sig0000039a,
      DI => blk00000003_sig0000039d,
      S => blk00000003_sig0000039b,
      O => blk00000003_sig0000038e
    );
  blk00000003_blk00000267 : XORCY
    port map (
      CI => blk00000003_sig0000039a,
      LI => blk00000003_sig0000039b,
      O => blk00000003_sig0000039c
    );
  blk00000003_blk00000266 : MUXCY
    port map (
      CI => blk00000003_sig00000379,
      DI => blk00000003_sig00000398,
      S => blk00000003_sig0000037a,
      O => blk00000003_sig00000399
    );
  blk00000003_blk00000265 : MUXCY
    port map (
      CI => blk00000003_sig0000038e,
      DI => blk00000003_sig00000397,
      S => blk00000003_sig0000038f,
      O => blk00000003_sig0000038b
    );
  blk00000003_blk00000264 : MUXCY
    port map (
      CI => blk00000003_sig0000038b,
      DI => blk00000003_sig00000396,
      S => blk00000003_sig0000038c,
      O => blk00000003_sig00000388
    );
  blk00000003_blk00000263 : MUXCY
    port map (
      CI => blk00000003_sig00000388,
      DI => blk00000003_sig00000395,
      S => blk00000003_sig00000389,
      O => blk00000003_sig00000385
    );
  blk00000003_blk00000262 : MUXCY
    port map (
      CI => blk00000003_sig00000385,
      DI => blk00000003_sig00000394,
      S => blk00000003_sig00000386,
      O => blk00000003_sig00000382
    );
  blk00000003_blk00000261 : MUXCY
    port map (
      CI => blk00000003_sig00000382,
      DI => blk00000003_sig00000393,
      S => blk00000003_sig00000383,
      O => blk00000003_sig0000037f
    );
  blk00000003_blk00000260 : MUXCY
    port map (
      CI => blk00000003_sig0000037f,
      DI => blk00000003_sig00000392,
      S => blk00000003_sig00000380,
      O => blk00000003_sig0000037c
    );
  blk00000003_blk0000025f : MUXCY
    port map (
      CI => blk00000003_sig0000037c,
      DI => blk00000003_sig00000391,
      S => blk00000003_sig0000037d,
      O => blk00000003_sig00000379
    );
  blk00000003_blk0000025e : XORCY
    port map (
      CI => blk00000003_sig0000038e,
      LI => blk00000003_sig0000038f,
      O => blk00000003_sig00000390
    );
  blk00000003_blk0000025d : XORCY
    port map (
      CI => blk00000003_sig0000038b,
      LI => blk00000003_sig0000038c,
      O => blk00000003_sig0000038d
    );
  blk00000003_blk0000025c : XORCY
    port map (
      CI => blk00000003_sig00000388,
      LI => blk00000003_sig00000389,
      O => blk00000003_sig0000038a
    );
  blk00000003_blk0000025b : XORCY
    port map (
      CI => blk00000003_sig00000385,
      LI => blk00000003_sig00000386,
      O => blk00000003_sig00000387
    );
  blk00000003_blk0000025a : XORCY
    port map (
      CI => blk00000003_sig00000382,
      LI => blk00000003_sig00000383,
      O => blk00000003_sig00000384
    );
  blk00000003_blk00000259 : XORCY
    port map (
      CI => blk00000003_sig0000037f,
      LI => blk00000003_sig00000380,
      O => blk00000003_sig00000381
    );
  blk00000003_blk00000258 : XORCY
    port map (
      CI => blk00000003_sig0000037c,
      LI => blk00000003_sig0000037d,
      O => blk00000003_sig0000037e
    );
  blk00000003_blk00000257 : XORCY
    port map (
      CI => blk00000003_sig00000379,
      LI => blk00000003_sig0000037a,
      O => blk00000003_sig0000037b
    );
  blk00000003_blk00000256 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000373,
      Q => blk00000003_sig00000378
    );
  blk00000003_blk00000255 : MUXCY
    port map (
      CI => blk00000003_sig00000374,
      DI => blk00000003_sig00000377,
      S => blk00000003_sig00000375,
      O => blk00000003_sig00000368
    );
  blk00000003_blk00000254 : XORCY
    port map (
      CI => blk00000003_sig00000374,
      LI => blk00000003_sig00000375,
      O => blk00000003_sig00000376
    );
  blk00000003_blk00000253 : MUXCY
    port map (
      CI => blk00000003_sig00000353,
      DI => blk00000003_sig00000372,
      S => blk00000003_sig00000354,
      O => blk00000003_sig00000373
    );
  blk00000003_blk00000252 : MUXCY
    port map (
      CI => blk00000003_sig00000368,
      DI => blk00000003_sig00000371,
      S => blk00000003_sig00000369,
      O => blk00000003_sig00000365
    );
  blk00000003_blk00000251 : MUXCY
    port map (
      CI => blk00000003_sig00000365,
      DI => blk00000003_sig00000370,
      S => blk00000003_sig00000366,
      O => blk00000003_sig00000362
    );
  blk00000003_blk00000250 : MUXCY
    port map (
      CI => blk00000003_sig00000362,
      DI => blk00000003_sig0000036f,
      S => blk00000003_sig00000363,
      O => blk00000003_sig0000035f
    );
  blk00000003_blk0000024f : MUXCY
    port map (
      CI => blk00000003_sig0000035f,
      DI => blk00000003_sig0000036e,
      S => blk00000003_sig00000360,
      O => blk00000003_sig0000035c
    );
  blk00000003_blk0000024e : MUXCY
    port map (
      CI => blk00000003_sig0000035c,
      DI => blk00000003_sig0000036d,
      S => blk00000003_sig0000035d,
      O => blk00000003_sig00000359
    );
  blk00000003_blk0000024d : MUXCY
    port map (
      CI => blk00000003_sig00000359,
      DI => blk00000003_sig0000036c,
      S => blk00000003_sig0000035a,
      O => blk00000003_sig00000356
    );
  blk00000003_blk0000024c : MUXCY
    port map (
      CI => blk00000003_sig00000356,
      DI => blk00000003_sig0000036b,
      S => blk00000003_sig00000357,
      O => blk00000003_sig00000353
    );
  blk00000003_blk0000024b : XORCY
    port map (
      CI => blk00000003_sig00000368,
      LI => blk00000003_sig00000369,
      O => blk00000003_sig0000036a
    );
  blk00000003_blk0000024a : XORCY
    port map (
      CI => blk00000003_sig00000365,
      LI => blk00000003_sig00000366,
      O => blk00000003_sig00000367
    );
  blk00000003_blk00000249 : XORCY
    port map (
      CI => blk00000003_sig00000362,
      LI => blk00000003_sig00000363,
      O => blk00000003_sig00000364
    );
  blk00000003_blk00000248 : XORCY
    port map (
      CI => blk00000003_sig0000035f,
      LI => blk00000003_sig00000360,
      O => blk00000003_sig00000361
    );
  blk00000003_blk00000247 : XORCY
    port map (
      CI => blk00000003_sig0000035c,
      LI => blk00000003_sig0000035d,
      O => blk00000003_sig0000035e
    );
  blk00000003_blk00000246 : XORCY
    port map (
      CI => blk00000003_sig00000359,
      LI => blk00000003_sig0000035a,
      O => blk00000003_sig0000035b
    );
  blk00000003_blk00000245 : XORCY
    port map (
      CI => blk00000003_sig00000356,
      LI => blk00000003_sig00000357,
      O => blk00000003_sig00000358
    );
  blk00000003_blk00000244 : XORCY
    port map (
      CI => blk00000003_sig00000353,
      LI => blk00000003_sig00000354,
      O => blk00000003_sig00000355
    );
  blk00000003_blk00000243 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000034d,
      Q => blk00000003_sig00000352
    );
  blk00000003_blk00000242 : MUXCY
    port map (
      CI => blk00000003_sig0000034e,
      DI => blk00000003_sig00000351,
      S => blk00000003_sig0000034f,
      O => blk00000003_sig00000342
    );
  blk00000003_blk00000241 : XORCY
    port map (
      CI => blk00000003_sig0000034e,
      LI => blk00000003_sig0000034f,
      O => blk00000003_sig00000350
    );
  blk00000003_blk00000240 : MUXCY
    port map (
      CI => blk00000003_sig0000032d,
      DI => blk00000003_sig0000034c,
      S => blk00000003_sig0000032e,
      O => blk00000003_sig0000034d
    );
  blk00000003_blk0000023f : MUXCY
    port map (
      CI => blk00000003_sig00000342,
      DI => blk00000003_sig0000034b,
      S => blk00000003_sig00000343,
      O => blk00000003_sig0000033f
    );
  blk00000003_blk0000023e : MUXCY
    port map (
      CI => blk00000003_sig0000033f,
      DI => blk00000003_sig0000034a,
      S => blk00000003_sig00000340,
      O => blk00000003_sig0000033c
    );
  blk00000003_blk0000023d : MUXCY
    port map (
      CI => blk00000003_sig0000033c,
      DI => blk00000003_sig00000349,
      S => blk00000003_sig0000033d,
      O => blk00000003_sig00000339
    );
  blk00000003_blk0000023c : MUXCY
    port map (
      CI => blk00000003_sig00000339,
      DI => blk00000003_sig00000348,
      S => blk00000003_sig0000033a,
      O => blk00000003_sig00000336
    );
  blk00000003_blk0000023b : MUXCY
    port map (
      CI => blk00000003_sig00000336,
      DI => blk00000003_sig00000347,
      S => blk00000003_sig00000337,
      O => blk00000003_sig00000333
    );
  blk00000003_blk0000023a : MUXCY
    port map (
      CI => blk00000003_sig00000333,
      DI => blk00000003_sig00000346,
      S => blk00000003_sig00000334,
      O => blk00000003_sig00000330
    );
  blk00000003_blk00000239 : MUXCY
    port map (
      CI => blk00000003_sig00000330,
      DI => blk00000003_sig00000345,
      S => blk00000003_sig00000331,
      O => blk00000003_sig0000032d
    );
  blk00000003_blk00000238 : XORCY
    port map (
      CI => blk00000003_sig00000342,
      LI => blk00000003_sig00000343,
      O => blk00000003_sig00000344
    );
  blk00000003_blk00000237 : XORCY
    port map (
      CI => blk00000003_sig0000033f,
      LI => blk00000003_sig00000340,
      O => blk00000003_sig00000341
    );
  blk00000003_blk00000236 : XORCY
    port map (
      CI => blk00000003_sig0000033c,
      LI => blk00000003_sig0000033d,
      O => blk00000003_sig0000033e
    );
  blk00000003_blk00000235 : XORCY
    port map (
      CI => blk00000003_sig00000339,
      LI => blk00000003_sig0000033a,
      O => blk00000003_sig0000033b
    );
  blk00000003_blk00000234 : XORCY
    port map (
      CI => blk00000003_sig00000336,
      LI => blk00000003_sig00000337,
      O => blk00000003_sig00000338
    );
  blk00000003_blk00000233 : XORCY
    port map (
      CI => blk00000003_sig00000333,
      LI => blk00000003_sig00000334,
      O => blk00000003_sig00000335
    );
  blk00000003_blk00000232 : XORCY
    port map (
      CI => blk00000003_sig00000330,
      LI => blk00000003_sig00000331,
      O => blk00000003_sig00000332
    );
  blk00000003_blk00000231 : XORCY
    port map (
      CI => blk00000003_sig0000032d,
      LI => blk00000003_sig0000032e,
      O => blk00000003_sig0000032f
    );
  blk00000003_blk00000230 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000327,
      Q => blk00000003_sig0000032c
    );
  blk00000003_blk0000022f : MUXCY
    port map (
      CI => blk00000003_sig00000328,
      DI => blk00000003_sig0000032b,
      S => blk00000003_sig00000329,
      O => blk00000003_sig0000031c
    );
  blk00000003_blk0000022e : XORCY
    port map (
      CI => blk00000003_sig00000328,
      LI => blk00000003_sig00000329,
      O => blk00000003_sig0000032a
    );
  blk00000003_blk0000022d : MUXCY
    port map (
      CI => blk00000003_sig00000307,
      DI => blk00000003_sig00000326,
      S => blk00000003_sig00000308,
      O => blk00000003_sig00000327
    );
  blk00000003_blk0000022c : MUXCY
    port map (
      CI => blk00000003_sig0000031c,
      DI => blk00000003_sig00000325,
      S => blk00000003_sig0000031d,
      O => blk00000003_sig00000319
    );
  blk00000003_blk0000022b : MUXCY
    port map (
      CI => blk00000003_sig00000319,
      DI => blk00000003_sig00000324,
      S => blk00000003_sig0000031a,
      O => blk00000003_sig00000316
    );
  blk00000003_blk0000022a : MUXCY
    port map (
      CI => blk00000003_sig00000316,
      DI => blk00000003_sig00000323,
      S => blk00000003_sig00000317,
      O => blk00000003_sig00000313
    );
  blk00000003_blk00000229 : MUXCY
    port map (
      CI => blk00000003_sig00000313,
      DI => blk00000003_sig00000322,
      S => blk00000003_sig00000314,
      O => blk00000003_sig00000310
    );
  blk00000003_blk00000228 : MUXCY
    port map (
      CI => blk00000003_sig00000310,
      DI => blk00000003_sig00000321,
      S => blk00000003_sig00000311,
      O => blk00000003_sig0000030d
    );
  blk00000003_blk00000227 : MUXCY
    port map (
      CI => blk00000003_sig0000030d,
      DI => blk00000003_sig00000320,
      S => blk00000003_sig0000030e,
      O => blk00000003_sig0000030a
    );
  blk00000003_blk00000226 : MUXCY
    port map (
      CI => blk00000003_sig0000030a,
      DI => blk00000003_sig0000031f,
      S => blk00000003_sig0000030b,
      O => blk00000003_sig00000307
    );
  blk00000003_blk00000225 : XORCY
    port map (
      CI => blk00000003_sig0000031c,
      LI => blk00000003_sig0000031d,
      O => blk00000003_sig0000031e
    );
  blk00000003_blk00000224 : XORCY
    port map (
      CI => blk00000003_sig00000319,
      LI => blk00000003_sig0000031a,
      O => blk00000003_sig0000031b
    );
  blk00000003_blk00000223 : XORCY
    port map (
      CI => blk00000003_sig00000316,
      LI => blk00000003_sig00000317,
      O => blk00000003_sig00000318
    );
  blk00000003_blk00000222 : XORCY
    port map (
      CI => blk00000003_sig00000313,
      LI => blk00000003_sig00000314,
      O => blk00000003_sig00000315
    );
  blk00000003_blk00000221 : XORCY
    port map (
      CI => blk00000003_sig00000310,
      LI => blk00000003_sig00000311,
      O => blk00000003_sig00000312
    );
  blk00000003_blk00000220 : XORCY
    port map (
      CI => blk00000003_sig0000030d,
      LI => blk00000003_sig0000030e,
      O => blk00000003_sig0000030f
    );
  blk00000003_blk0000021f : XORCY
    port map (
      CI => blk00000003_sig0000030a,
      LI => blk00000003_sig0000030b,
      O => blk00000003_sig0000030c
    );
  blk00000003_blk0000021e : XORCY
    port map (
      CI => blk00000003_sig00000307,
      LI => blk00000003_sig00000308,
      O => blk00000003_sig00000309
    );
  blk00000003_blk0000021d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000301,
      Q => blk00000003_sig00000306
    );
  blk00000003_blk0000021c : MUXCY
    port map (
      CI => blk00000003_sig00000302,
      DI => blk00000003_sig00000305,
      S => blk00000003_sig00000303,
      O => blk00000003_sig000002f6
    );
  blk00000003_blk0000021b : XORCY
    port map (
      CI => blk00000003_sig00000302,
      LI => blk00000003_sig00000303,
      O => blk00000003_sig00000304
    );
  blk00000003_blk0000021a : MUXCY
    port map (
      CI => blk00000003_sig000002e1,
      DI => blk00000003_sig00000300,
      S => blk00000003_sig000002e2,
      O => blk00000003_sig00000301
    );
  blk00000003_blk00000219 : MUXCY
    port map (
      CI => blk00000003_sig000002f6,
      DI => blk00000003_sig000002ff,
      S => blk00000003_sig000002f7,
      O => blk00000003_sig000002f3
    );
  blk00000003_blk00000218 : MUXCY
    port map (
      CI => blk00000003_sig000002f3,
      DI => blk00000003_sig000002fe,
      S => blk00000003_sig000002f4,
      O => blk00000003_sig000002f0
    );
  blk00000003_blk00000217 : MUXCY
    port map (
      CI => blk00000003_sig000002f0,
      DI => blk00000003_sig000002fd,
      S => blk00000003_sig000002f1,
      O => blk00000003_sig000002ed
    );
  blk00000003_blk00000216 : MUXCY
    port map (
      CI => blk00000003_sig000002ed,
      DI => blk00000003_sig000002fc,
      S => blk00000003_sig000002ee,
      O => blk00000003_sig000002ea
    );
  blk00000003_blk00000215 : MUXCY
    port map (
      CI => blk00000003_sig000002ea,
      DI => blk00000003_sig000002fb,
      S => blk00000003_sig000002eb,
      O => blk00000003_sig000002e7
    );
  blk00000003_blk00000214 : MUXCY
    port map (
      CI => blk00000003_sig000002e7,
      DI => blk00000003_sig000002fa,
      S => blk00000003_sig000002e8,
      O => blk00000003_sig000002e4
    );
  blk00000003_blk00000213 : MUXCY
    port map (
      CI => blk00000003_sig000002e4,
      DI => blk00000003_sig000002f9,
      S => blk00000003_sig000002e5,
      O => blk00000003_sig000002e1
    );
  blk00000003_blk00000212 : XORCY
    port map (
      CI => blk00000003_sig000002f6,
      LI => blk00000003_sig000002f7,
      O => blk00000003_sig000002f8
    );
  blk00000003_blk00000211 : XORCY
    port map (
      CI => blk00000003_sig000002f3,
      LI => blk00000003_sig000002f4,
      O => blk00000003_sig000002f5
    );
  blk00000003_blk00000210 : XORCY
    port map (
      CI => blk00000003_sig000002f0,
      LI => blk00000003_sig000002f1,
      O => blk00000003_sig000002f2
    );
  blk00000003_blk0000020f : XORCY
    port map (
      CI => blk00000003_sig000002ed,
      LI => blk00000003_sig000002ee,
      O => blk00000003_sig000002ef
    );
  blk00000003_blk0000020e : XORCY
    port map (
      CI => blk00000003_sig000002ea,
      LI => blk00000003_sig000002eb,
      O => blk00000003_sig000002ec
    );
  blk00000003_blk0000020d : XORCY
    port map (
      CI => blk00000003_sig000002e7,
      LI => blk00000003_sig000002e8,
      O => blk00000003_sig000002e9
    );
  blk00000003_blk0000020c : XORCY
    port map (
      CI => blk00000003_sig000002e4,
      LI => blk00000003_sig000002e5,
      O => blk00000003_sig000002e6
    );
  blk00000003_blk0000020b : XORCY
    port map (
      CI => blk00000003_sig000002e1,
      LI => blk00000003_sig000002e2,
      O => blk00000003_sig000002e3
    );
  blk00000003_blk0000020a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002db,
      Q => blk00000003_sig000002e0
    );
  blk00000003_blk00000209 : MUXCY
    port map (
      CI => blk00000003_sig000002dc,
      DI => blk00000003_sig000002df,
      S => blk00000003_sig000002dd,
      O => blk00000003_sig000002d0
    );
  blk00000003_blk00000208 : XORCY
    port map (
      CI => blk00000003_sig000002dc,
      LI => blk00000003_sig000002dd,
      O => blk00000003_sig000002de
    );
  blk00000003_blk00000207 : MUXCY
    port map (
      CI => blk00000003_sig000002bb,
      DI => blk00000003_sig000002da,
      S => blk00000003_sig000002bc,
      O => blk00000003_sig000002db
    );
  blk00000003_blk00000206 : MUXCY
    port map (
      CI => blk00000003_sig000002d0,
      DI => blk00000003_sig000002d9,
      S => blk00000003_sig000002d1,
      O => blk00000003_sig000002cd
    );
  blk00000003_blk00000205 : MUXCY
    port map (
      CI => blk00000003_sig000002cd,
      DI => blk00000003_sig000002d8,
      S => blk00000003_sig000002ce,
      O => blk00000003_sig000002ca
    );
  blk00000003_blk00000204 : MUXCY
    port map (
      CI => blk00000003_sig000002ca,
      DI => blk00000003_sig000002d7,
      S => blk00000003_sig000002cb,
      O => blk00000003_sig000002c7
    );
  blk00000003_blk00000203 : MUXCY
    port map (
      CI => blk00000003_sig000002c7,
      DI => blk00000003_sig000002d6,
      S => blk00000003_sig000002c8,
      O => blk00000003_sig000002c4
    );
  blk00000003_blk00000202 : MUXCY
    port map (
      CI => blk00000003_sig000002c4,
      DI => blk00000003_sig000002d5,
      S => blk00000003_sig000002c5,
      O => blk00000003_sig000002c1
    );
  blk00000003_blk00000201 : MUXCY
    port map (
      CI => blk00000003_sig000002c1,
      DI => blk00000003_sig000002d4,
      S => blk00000003_sig000002c2,
      O => blk00000003_sig000002be
    );
  blk00000003_blk00000200 : MUXCY
    port map (
      CI => blk00000003_sig000002be,
      DI => blk00000003_sig000002d3,
      S => blk00000003_sig000002bf,
      O => blk00000003_sig000002bb
    );
  blk00000003_blk000001ff : XORCY
    port map (
      CI => blk00000003_sig000002d0,
      LI => blk00000003_sig000002d1,
      O => blk00000003_sig000002d2
    );
  blk00000003_blk000001fe : XORCY
    port map (
      CI => blk00000003_sig000002cd,
      LI => blk00000003_sig000002ce,
      O => blk00000003_sig000002cf
    );
  blk00000003_blk000001fd : XORCY
    port map (
      CI => blk00000003_sig000002ca,
      LI => blk00000003_sig000002cb,
      O => blk00000003_sig000002cc
    );
  blk00000003_blk000001fc : XORCY
    port map (
      CI => blk00000003_sig000002c7,
      LI => blk00000003_sig000002c8,
      O => blk00000003_sig000002c9
    );
  blk00000003_blk000001fb : XORCY
    port map (
      CI => blk00000003_sig000002c4,
      LI => blk00000003_sig000002c5,
      O => blk00000003_sig000002c6
    );
  blk00000003_blk000001fa : XORCY
    port map (
      CI => blk00000003_sig000002c1,
      LI => blk00000003_sig000002c2,
      O => blk00000003_sig000002c3
    );
  blk00000003_blk000001f9 : XORCY
    port map (
      CI => blk00000003_sig000002be,
      LI => blk00000003_sig000002bf,
      O => blk00000003_sig000002c0
    );
  blk00000003_blk000001f8 : XORCY
    port map (
      CI => blk00000003_sig000002bb,
      LI => blk00000003_sig000002bc,
      O => blk00000003_sig000002bd
    );
  blk00000003_blk000001f7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002b5,
      Q => blk00000003_sig000002ba
    );
  blk00000003_blk000001f6 : MUXCY
    port map (
      CI => blk00000003_sig000002b6,
      DI => blk00000003_sig000002b9,
      S => blk00000003_sig000002b7,
      O => blk00000003_sig000002aa
    );
  blk00000003_blk000001f5 : XORCY
    port map (
      CI => blk00000003_sig000002b6,
      LI => blk00000003_sig000002b7,
      O => blk00000003_sig000002b8
    );
  blk00000003_blk000001f4 : MUXCY
    port map (
      CI => blk00000003_sig00000295,
      DI => blk00000003_sig000002b4,
      S => blk00000003_sig00000296,
      O => blk00000003_sig000002b5
    );
  blk00000003_blk000001f3 : MUXCY
    port map (
      CI => blk00000003_sig000002aa,
      DI => blk00000003_sig000002b3,
      S => blk00000003_sig000002ab,
      O => blk00000003_sig000002a7
    );
  blk00000003_blk000001f2 : MUXCY
    port map (
      CI => blk00000003_sig000002a7,
      DI => blk00000003_sig000002b2,
      S => blk00000003_sig000002a8,
      O => blk00000003_sig000002a4
    );
  blk00000003_blk000001f1 : MUXCY
    port map (
      CI => blk00000003_sig000002a4,
      DI => blk00000003_sig000002b1,
      S => blk00000003_sig000002a5,
      O => blk00000003_sig000002a1
    );
  blk00000003_blk000001f0 : MUXCY
    port map (
      CI => blk00000003_sig000002a1,
      DI => blk00000003_sig000002b0,
      S => blk00000003_sig000002a2,
      O => blk00000003_sig0000029e
    );
  blk00000003_blk000001ef : MUXCY
    port map (
      CI => blk00000003_sig0000029e,
      DI => blk00000003_sig000002af,
      S => blk00000003_sig0000029f,
      O => blk00000003_sig0000029b
    );
  blk00000003_blk000001ee : MUXCY
    port map (
      CI => blk00000003_sig0000029b,
      DI => blk00000003_sig000002ae,
      S => blk00000003_sig0000029c,
      O => blk00000003_sig00000298
    );
  blk00000003_blk000001ed : MUXCY
    port map (
      CI => blk00000003_sig00000298,
      DI => blk00000003_sig000002ad,
      S => blk00000003_sig00000299,
      O => blk00000003_sig00000295
    );
  blk00000003_blk000001ec : XORCY
    port map (
      CI => blk00000003_sig000002aa,
      LI => blk00000003_sig000002ab,
      O => blk00000003_sig000002ac
    );
  blk00000003_blk000001eb : XORCY
    port map (
      CI => blk00000003_sig000002a7,
      LI => blk00000003_sig000002a8,
      O => blk00000003_sig000002a9
    );
  blk00000003_blk000001ea : XORCY
    port map (
      CI => blk00000003_sig000002a4,
      LI => blk00000003_sig000002a5,
      O => blk00000003_sig000002a6
    );
  blk00000003_blk000001e9 : XORCY
    port map (
      CI => blk00000003_sig000002a1,
      LI => blk00000003_sig000002a2,
      O => blk00000003_sig000002a3
    );
  blk00000003_blk000001e8 : XORCY
    port map (
      CI => blk00000003_sig0000029e,
      LI => blk00000003_sig0000029f,
      O => blk00000003_sig000002a0
    );
  blk00000003_blk000001e7 : XORCY
    port map (
      CI => blk00000003_sig0000029b,
      LI => blk00000003_sig0000029c,
      O => blk00000003_sig0000029d
    );
  blk00000003_blk000001e6 : XORCY
    port map (
      CI => blk00000003_sig00000298,
      LI => blk00000003_sig00000299,
      O => blk00000003_sig0000029a
    );
  blk00000003_blk000001e5 : XORCY
    port map (
      CI => blk00000003_sig00000295,
      LI => blk00000003_sig00000296,
      O => blk00000003_sig00000297
    );
  blk00000003_blk000001e4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000028f,
      Q => blk00000003_sig00000294
    );
  blk00000003_blk000001e3 : MUXCY
    port map (
      CI => blk00000003_sig00000290,
      DI => blk00000003_sig00000293,
      S => blk00000003_sig00000291,
      O => blk00000003_sig00000284
    );
  blk00000003_blk000001e2 : XORCY
    port map (
      CI => blk00000003_sig00000290,
      LI => blk00000003_sig00000291,
      O => blk00000003_sig00000292
    );
  blk00000003_blk000001e1 : MUXCY
    port map (
      CI => blk00000003_sig0000026f,
      DI => blk00000003_sig0000028e,
      S => blk00000003_sig00000270,
      O => blk00000003_sig0000028f
    );
  blk00000003_blk000001e0 : MUXCY
    port map (
      CI => blk00000003_sig00000284,
      DI => blk00000003_sig0000028d,
      S => blk00000003_sig00000285,
      O => blk00000003_sig00000281
    );
  blk00000003_blk000001df : MUXCY
    port map (
      CI => blk00000003_sig00000281,
      DI => blk00000003_sig0000028c,
      S => blk00000003_sig00000282,
      O => blk00000003_sig0000027e
    );
  blk00000003_blk000001de : MUXCY
    port map (
      CI => blk00000003_sig0000027e,
      DI => blk00000003_sig0000028b,
      S => blk00000003_sig0000027f,
      O => blk00000003_sig0000027b
    );
  blk00000003_blk000001dd : MUXCY
    port map (
      CI => blk00000003_sig0000027b,
      DI => blk00000003_sig0000028a,
      S => blk00000003_sig0000027c,
      O => blk00000003_sig00000278
    );
  blk00000003_blk000001dc : MUXCY
    port map (
      CI => blk00000003_sig00000278,
      DI => blk00000003_sig00000289,
      S => blk00000003_sig00000279,
      O => blk00000003_sig00000275
    );
  blk00000003_blk000001db : MUXCY
    port map (
      CI => blk00000003_sig00000275,
      DI => blk00000003_sig00000288,
      S => blk00000003_sig00000276,
      O => blk00000003_sig00000272
    );
  blk00000003_blk000001da : MUXCY
    port map (
      CI => blk00000003_sig00000272,
      DI => blk00000003_sig00000287,
      S => blk00000003_sig00000273,
      O => blk00000003_sig0000026f
    );
  blk00000003_blk000001d9 : XORCY
    port map (
      CI => blk00000003_sig00000284,
      LI => blk00000003_sig00000285,
      O => blk00000003_sig00000286
    );
  blk00000003_blk000001d8 : XORCY
    port map (
      CI => blk00000003_sig00000281,
      LI => blk00000003_sig00000282,
      O => blk00000003_sig00000283
    );
  blk00000003_blk000001d7 : XORCY
    port map (
      CI => blk00000003_sig0000027e,
      LI => blk00000003_sig0000027f,
      O => blk00000003_sig00000280
    );
  blk00000003_blk000001d6 : XORCY
    port map (
      CI => blk00000003_sig0000027b,
      LI => blk00000003_sig0000027c,
      O => blk00000003_sig0000027d
    );
  blk00000003_blk000001d5 : XORCY
    port map (
      CI => blk00000003_sig00000278,
      LI => blk00000003_sig00000279,
      O => blk00000003_sig0000027a
    );
  blk00000003_blk000001d4 : XORCY
    port map (
      CI => blk00000003_sig00000275,
      LI => blk00000003_sig00000276,
      O => blk00000003_sig00000277
    );
  blk00000003_blk000001d3 : XORCY
    port map (
      CI => blk00000003_sig00000272,
      LI => blk00000003_sig00000273,
      O => blk00000003_sig00000274
    );
  blk00000003_blk000001d2 : XORCY
    port map (
      CI => blk00000003_sig0000026f,
      LI => blk00000003_sig00000270,
      O => blk00000003_sig00000271
    );
  blk00000003_blk000001d1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000269,
      Q => blk00000003_sig0000026e
    );
  blk00000003_blk000001d0 : MUXCY
    port map (
      CI => blk00000003_sig0000026a,
      DI => blk00000003_sig0000026d,
      S => blk00000003_sig0000026b,
      O => blk00000003_sig0000025e
    );
  blk00000003_blk000001cf : XORCY
    port map (
      CI => blk00000003_sig0000026a,
      LI => blk00000003_sig0000026b,
      O => blk00000003_sig0000026c
    );
  blk00000003_blk000001ce : MUXCY
    port map (
      CI => blk00000003_sig00000249,
      DI => blk00000003_sig00000268,
      S => blk00000003_sig0000024a,
      O => blk00000003_sig00000269
    );
  blk00000003_blk000001cd : MUXCY
    port map (
      CI => blk00000003_sig0000025e,
      DI => blk00000003_sig00000267,
      S => blk00000003_sig0000025f,
      O => blk00000003_sig0000025b
    );
  blk00000003_blk000001cc : MUXCY
    port map (
      CI => blk00000003_sig0000025b,
      DI => blk00000003_sig00000266,
      S => blk00000003_sig0000025c,
      O => blk00000003_sig00000258
    );
  blk00000003_blk000001cb : MUXCY
    port map (
      CI => blk00000003_sig00000258,
      DI => blk00000003_sig00000265,
      S => blk00000003_sig00000259,
      O => blk00000003_sig00000255
    );
  blk00000003_blk000001ca : MUXCY
    port map (
      CI => blk00000003_sig00000255,
      DI => blk00000003_sig00000264,
      S => blk00000003_sig00000256,
      O => blk00000003_sig00000252
    );
  blk00000003_blk000001c9 : MUXCY
    port map (
      CI => blk00000003_sig00000252,
      DI => blk00000003_sig00000263,
      S => blk00000003_sig00000253,
      O => blk00000003_sig0000024f
    );
  blk00000003_blk000001c8 : MUXCY
    port map (
      CI => blk00000003_sig0000024f,
      DI => blk00000003_sig00000262,
      S => blk00000003_sig00000250,
      O => blk00000003_sig0000024c
    );
  blk00000003_blk000001c7 : MUXCY
    port map (
      CI => blk00000003_sig0000024c,
      DI => blk00000003_sig00000261,
      S => blk00000003_sig0000024d,
      O => blk00000003_sig00000249
    );
  blk00000003_blk000001c6 : XORCY
    port map (
      CI => blk00000003_sig0000025e,
      LI => blk00000003_sig0000025f,
      O => blk00000003_sig00000260
    );
  blk00000003_blk000001c5 : XORCY
    port map (
      CI => blk00000003_sig0000025b,
      LI => blk00000003_sig0000025c,
      O => blk00000003_sig0000025d
    );
  blk00000003_blk000001c4 : XORCY
    port map (
      CI => blk00000003_sig00000258,
      LI => blk00000003_sig00000259,
      O => blk00000003_sig0000025a
    );
  blk00000003_blk000001c3 : XORCY
    port map (
      CI => blk00000003_sig00000255,
      LI => blk00000003_sig00000256,
      O => blk00000003_sig00000257
    );
  blk00000003_blk000001c2 : XORCY
    port map (
      CI => blk00000003_sig00000252,
      LI => blk00000003_sig00000253,
      O => blk00000003_sig00000254
    );
  blk00000003_blk000001c1 : XORCY
    port map (
      CI => blk00000003_sig0000024f,
      LI => blk00000003_sig00000250,
      O => blk00000003_sig00000251
    );
  blk00000003_blk000001c0 : XORCY
    port map (
      CI => blk00000003_sig0000024c,
      LI => blk00000003_sig0000024d,
      O => blk00000003_sig0000024e
    );
  blk00000003_blk000001bf : XORCY
    port map (
      CI => blk00000003_sig00000249,
      LI => blk00000003_sig0000024a,
      O => blk00000003_sig0000024b
    );
  blk00000003_blk000001be : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000243,
      Q => blk00000003_sig00000248
    );
  blk00000003_blk000001bd : MUXCY
    port map (
      CI => blk00000003_sig00000244,
      DI => blk00000003_sig00000247,
      S => blk00000003_sig00000245,
      O => blk00000003_sig00000238
    );
  blk00000003_blk000001bc : XORCY
    port map (
      CI => blk00000003_sig00000244,
      LI => blk00000003_sig00000245,
      O => blk00000003_sig00000246
    );
  blk00000003_blk000001bb : MUXCY
    port map (
      CI => blk00000003_sig00000223,
      DI => blk00000003_sig00000242,
      S => blk00000003_sig00000224,
      O => blk00000003_sig00000243
    );
  blk00000003_blk000001ba : MUXCY
    port map (
      CI => blk00000003_sig00000238,
      DI => blk00000003_sig00000241,
      S => blk00000003_sig00000239,
      O => blk00000003_sig00000235
    );
  blk00000003_blk000001b9 : MUXCY
    port map (
      CI => blk00000003_sig00000235,
      DI => blk00000003_sig00000240,
      S => blk00000003_sig00000236,
      O => blk00000003_sig00000232
    );
  blk00000003_blk000001b8 : MUXCY
    port map (
      CI => blk00000003_sig00000232,
      DI => blk00000003_sig0000023f,
      S => blk00000003_sig00000233,
      O => blk00000003_sig0000022f
    );
  blk00000003_blk000001b7 : MUXCY
    port map (
      CI => blk00000003_sig0000022f,
      DI => blk00000003_sig0000023e,
      S => blk00000003_sig00000230,
      O => blk00000003_sig0000022c
    );
  blk00000003_blk000001b6 : MUXCY
    port map (
      CI => blk00000003_sig0000022c,
      DI => blk00000003_sig0000023d,
      S => blk00000003_sig0000022d,
      O => blk00000003_sig00000229
    );
  blk00000003_blk000001b5 : MUXCY
    port map (
      CI => blk00000003_sig00000229,
      DI => blk00000003_sig0000023c,
      S => blk00000003_sig0000022a,
      O => blk00000003_sig00000226
    );
  blk00000003_blk000001b4 : MUXCY
    port map (
      CI => blk00000003_sig00000226,
      DI => blk00000003_sig0000023b,
      S => blk00000003_sig00000227,
      O => blk00000003_sig00000223
    );
  blk00000003_blk000001b3 : XORCY
    port map (
      CI => blk00000003_sig00000238,
      LI => blk00000003_sig00000239,
      O => blk00000003_sig0000023a
    );
  blk00000003_blk000001b2 : XORCY
    port map (
      CI => blk00000003_sig00000235,
      LI => blk00000003_sig00000236,
      O => blk00000003_sig00000237
    );
  blk00000003_blk000001b1 : XORCY
    port map (
      CI => blk00000003_sig00000232,
      LI => blk00000003_sig00000233,
      O => blk00000003_sig00000234
    );
  blk00000003_blk000001b0 : XORCY
    port map (
      CI => blk00000003_sig0000022f,
      LI => blk00000003_sig00000230,
      O => blk00000003_sig00000231
    );
  blk00000003_blk000001af : XORCY
    port map (
      CI => blk00000003_sig0000022c,
      LI => blk00000003_sig0000022d,
      O => blk00000003_sig0000022e
    );
  blk00000003_blk000001ae : XORCY
    port map (
      CI => blk00000003_sig00000229,
      LI => blk00000003_sig0000022a,
      O => blk00000003_sig0000022b
    );
  blk00000003_blk000001ad : XORCY
    port map (
      CI => blk00000003_sig00000226,
      LI => blk00000003_sig00000227,
      O => blk00000003_sig00000228
    );
  blk00000003_blk000001ac : XORCY
    port map (
      CI => blk00000003_sig00000223,
      LI => blk00000003_sig00000224,
      O => blk00000003_sig00000225
    );
  blk00000003_blk000001ab : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000021d,
      Q => blk00000003_sig00000222
    );
  blk00000003_blk000001aa : MUXCY
    port map (
      CI => blk00000003_sig0000021e,
      DI => blk00000003_sig00000221,
      S => blk00000003_sig0000021f,
      O => blk00000003_sig00000212
    );
  blk00000003_blk000001a9 : XORCY
    port map (
      CI => blk00000003_sig0000021e,
      LI => blk00000003_sig0000021f,
      O => blk00000003_sig00000220
    );
  blk00000003_blk000001a8 : MUXCY
    port map (
      CI => blk00000003_sig000001fd,
      DI => blk00000003_sig0000021c,
      S => blk00000003_sig000001fe,
      O => blk00000003_sig0000021d
    );
  blk00000003_blk000001a7 : MUXCY
    port map (
      CI => blk00000003_sig00000212,
      DI => blk00000003_sig0000021b,
      S => blk00000003_sig00000213,
      O => blk00000003_sig0000020f
    );
  blk00000003_blk000001a6 : MUXCY
    port map (
      CI => blk00000003_sig0000020f,
      DI => blk00000003_sig0000021a,
      S => blk00000003_sig00000210,
      O => blk00000003_sig0000020c
    );
  blk00000003_blk000001a5 : MUXCY
    port map (
      CI => blk00000003_sig0000020c,
      DI => blk00000003_sig00000219,
      S => blk00000003_sig0000020d,
      O => blk00000003_sig00000209
    );
  blk00000003_blk000001a4 : MUXCY
    port map (
      CI => blk00000003_sig00000209,
      DI => blk00000003_sig00000218,
      S => blk00000003_sig0000020a,
      O => blk00000003_sig00000206
    );
  blk00000003_blk000001a3 : MUXCY
    port map (
      CI => blk00000003_sig00000206,
      DI => blk00000003_sig00000217,
      S => blk00000003_sig00000207,
      O => blk00000003_sig00000203
    );
  blk00000003_blk000001a2 : MUXCY
    port map (
      CI => blk00000003_sig00000203,
      DI => blk00000003_sig00000216,
      S => blk00000003_sig00000204,
      O => blk00000003_sig00000200
    );
  blk00000003_blk000001a1 : MUXCY
    port map (
      CI => blk00000003_sig00000200,
      DI => blk00000003_sig00000215,
      S => blk00000003_sig00000201,
      O => blk00000003_sig000001fd
    );
  blk00000003_blk000001a0 : XORCY
    port map (
      CI => blk00000003_sig00000212,
      LI => blk00000003_sig00000213,
      O => blk00000003_sig00000214
    );
  blk00000003_blk0000019f : XORCY
    port map (
      CI => blk00000003_sig0000020f,
      LI => blk00000003_sig00000210,
      O => blk00000003_sig00000211
    );
  blk00000003_blk0000019e : XORCY
    port map (
      CI => blk00000003_sig0000020c,
      LI => blk00000003_sig0000020d,
      O => blk00000003_sig0000020e
    );
  blk00000003_blk0000019d : XORCY
    port map (
      CI => blk00000003_sig00000209,
      LI => blk00000003_sig0000020a,
      O => blk00000003_sig0000020b
    );
  blk00000003_blk0000019c : XORCY
    port map (
      CI => blk00000003_sig00000206,
      LI => blk00000003_sig00000207,
      O => blk00000003_sig00000208
    );
  blk00000003_blk0000019b : XORCY
    port map (
      CI => blk00000003_sig00000203,
      LI => blk00000003_sig00000204,
      O => blk00000003_sig00000205
    );
  blk00000003_blk0000019a : XORCY
    port map (
      CI => blk00000003_sig00000200,
      LI => blk00000003_sig00000201,
      O => blk00000003_sig00000202
    );
  blk00000003_blk00000199 : XORCY
    port map (
      CI => blk00000003_sig000001fd,
      LI => blk00000003_sig000001fe,
      O => blk00000003_sig000001ff
    );
  blk00000003_blk00000198 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001f9,
      Q => blk00000003_sig000001fc
    );
  blk00000003_blk00000197 : MUXCY
    port map (
      CI => NlwRenamedSig_OI_rfd,
      DI => blk00000003_sig000000bb,
      S => blk00000003_sig000001fa,
      O => blk00000003_sig000001f6
    );
  blk00000003_blk00000196 : XORCY
    port map (
      CI => NlwRenamedSig_OI_rfd,
      LI => blk00000003_sig000001fa,
      O => blk00000003_sig000001fb
    );
  blk00000003_blk00000195 : MUXCY
    port map (
      CI => blk00000003_sig000001e3,
      DI => blk00000003_sig00000053,
      S => NlwRenamedSig_OI_rfd,
      O => blk00000003_sig000001f9
    );
  blk00000003_blk00000194 : MUXCY
    port map (
      CI => blk00000003_sig000001f6,
      DI => blk00000003_sig00000053,
      S => blk00000003_sig000001f7,
      O => blk00000003_sig000001f3
    );
  blk00000003_blk00000193 : MUXCY
    port map (
      CI => blk00000003_sig000001f3,
      DI => blk00000003_sig00000053,
      S => blk00000003_sig000001f4,
      O => blk00000003_sig000001f0
    );
  blk00000003_blk00000192 : MUXCY
    port map (
      CI => blk00000003_sig000001f0,
      DI => blk00000003_sig00000053,
      S => blk00000003_sig000001f1,
      O => blk00000003_sig000001ed
    );
  blk00000003_blk00000191 : MUXCY
    port map (
      CI => blk00000003_sig000001ed,
      DI => blk00000003_sig00000053,
      S => blk00000003_sig000001ee,
      O => blk00000003_sig000001ea
    );
  blk00000003_blk00000190 : MUXCY
    port map (
      CI => blk00000003_sig000001ea,
      DI => blk00000003_sig00000053,
      S => blk00000003_sig000001eb,
      O => blk00000003_sig000001e7
    );
  blk00000003_blk0000018f : MUXCY
    port map (
      CI => blk00000003_sig000001e7,
      DI => blk00000003_sig00000053,
      S => blk00000003_sig000001e8,
      O => blk00000003_sig000001e4
    );
  blk00000003_blk0000018e : MUXCY
    port map (
      CI => blk00000003_sig000001e4,
      DI => blk00000003_sig00000053,
      S => blk00000003_sig000001e5,
      O => blk00000003_sig000001e3
    );
  blk00000003_blk0000018d : XORCY
    port map (
      CI => blk00000003_sig000001f6,
      LI => blk00000003_sig000001f7,
      O => blk00000003_sig000001f8
    );
  blk00000003_blk0000018c : XORCY
    port map (
      CI => blk00000003_sig000001f3,
      LI => blk00000003_sig000001f4,
      O => blk00000003_sig000001f5
    );
  blk00000003_blk0000018b : XORCY
    port map (
      CI => blk00000003_sig000001f0,
      LI => blk00000003_sig000001f1,
      O => blk00000003_sig000001f2
    );
  blk00000003_blk0000018a : XORCY
    port map (
      CI => blk00000003_sig000001ed,
      LI => blk00000003_sig000001ee,
      O => blk00000003_sig000001ef
    );
  blk00000003_blk00000189 : XORCY
    port map (
      CI => blk00000003_sig000001ea,
      LI => blk00000003_sig000001eb,
      O => blk00000003_sig000001ec
    );
  blk00000003_blk00000188 : XORCY
    port map (
      CI => blk00000003_sig000001e7,
      LI => blk00000003_sig000001e8,
      O => blk00000003_sig000001e9
    );
  blk00000003_blk00000187 : XORCY
    port map (
      CI => blk00000003_sig000001e4,
      LI => blk00000003_sig000001e5,
      O => blk00000003_sig000001e6
    );
  blk00000003_blk00000186 : XORCY
    port map (
      CI => blk00000003_sig000001e3,
      LI => NlwRenamedSig_OI_rfd,
      O => NLW_blk00000003_blk00000186_O_UNCONNECTED
    );
  blk00000003_blk00000185 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(0),
      Q => blk00000003_sig000001e2
    );
  blk00000003_blk00000184 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(1),
      Q => blk00000003_sig000001e1
    );
  blk00000003_blk00000183 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(2),
      Q => blk00000003_sig000001e0
    );
  blk00000003_blk00000182 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(3),
      Q => blk00000003_sig000001df
    );
  blk00000003_blk00000181 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(4),
      Q => blk00000003_sig000001de
    );
  blk00000003_blk00000180 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(5),
      Q => blk00000003_sig000001dd
    );
  blk00000003_blk0000017f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(6),
      Q => blk00000003_sig000001dc
    );
  blk00000003_blk0000017e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(7),
      Q => blk00000003_sig000001db
    );
  blk00000003_blk0000017d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001e2,
      Q => blk00000003_sig000001da
    );
  blk00000003_blk0000017c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001e1,
      Q => blk00000003_sig000001d9
    );
  blk00000003_blk0000017b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001e0,
      Q => blk00000003_sig000001d8
    );
  blk00000003_blk0000017a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001df,
      Q => blk00000003_sig000001d7
    );
  blk00000003_blk00000179 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001de,
      Q => blk00000003_sig000001d6
    );
  blk00000003_blk00000178 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001dd,
      Q => blk00000003_sig000001d5
    );
  blk00000003_blk00000177 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001dc,
      Q => blk00000003_sig000001d4
    );
  blk00000003_blk00000176 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001db,
      Q => blk00000003_sig000001d3
    );
  blk00000003_blk00000175 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001da,
      Q => blk00000003_sig000001d2
    );
  blk00000003_blk00000174 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001d9,
      Q => blk00000003_sig000001d1
    );
  blk00000003_blk00000173 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001d8,
      Q => blk00000003_sig000001d0
    );
  blk00000003_blk00000172 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001d7,
      Q => blk00000003_sig000001cf
    );
  blk00000003_blk00000171 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001d6,
      Q => blk00000003_sig000001ce
    );
  blk00000003_blk00000170 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001d5,
      Q => blk00000003_sig000001cd
    );
  blk00000003_blk0000016f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001d4,
      Q => blk00000003_sig000001cc
    );
  blk00000003_blk0000016e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001d3,
      Q => blk00000003_sig000001cb
    );
  blk00000003_blk0000016d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001d2,
      Q => blk00000003_sig000001ca
    );
  blk00000003_blk0000016c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001d1,
      Q => blk00000003_sig000001c9
    );
  blk00000003_blk0000016b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001d0,
      Q => blk00000003_sig000001c8
    );
  blk00000003_blk0000016a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001cf,
      Q => blk00000003_sig000001c7
    );
  blk00000003_blk00000169 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001ce,
      Q => blk00000003_sig000001c6
    );
  blk00000003_blk00000168 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001cd,
      Q => blk00000003_sig000001c5
    );
  blk00000003_blk00000167 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001cc,
      Q => blk00000003_sig000001c4
    );
  blk00000003_blk00000166 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001cb,
      Q => blk00000003_sig000001c3
    );
  blk00000003_blk00000165 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001ca,
      Q => blk00000003_sig000001c2
    );
  blk00000003_blk00000164 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001c9,
      Q => blk00000003_sig000001c1
    );
  blk00000003_blk00000163 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001c8,
      Q => blk00000003_sig000001c0
    );
  blk00000003_blk00000162 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001c7,
      Q => blk00000003_sig000001bf
    );
  blk00000003_blk00000161 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001c6,
      Q => blk00000003_sig000001be
    );
  blk00000003_blk00000160 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001c5,
      Q => blk00000003_sig000001bd
    );
  blk00000003_blk0000015f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001c4,
      Q => blk00000003_sig000001bc
    );
  blk00000003_blk0000015e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001c3,
      Q => blk00000003_sig000001bb
    );
  blk00000003_blk0000015d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001c2,
      Q => blk00000003_sig000001ba
    );
  blk00000003_blk0000015c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001c1,
      Q => blk00000003_sig000001b9
    );
  blk00000003_blk0000015b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001c0,
      Q => blk00000003_sig000001b8
    );
  blk00000003_blk0000015a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001bf,
      Q => blk00000003_sig000001b7
    );
  blk00000003_blk00000159 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001be,
      Q => blk00000003_sig000001b6
    );
  blk00000003_blk00000158 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001bd,
      Q => blk00000003_sig000001b5
    );
  blk00000003_blk00000157 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001bc,
      Q => blk00000003_sig000001b4
    );
  blk00000003_blk00000156 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001bb,
      Q => blk00000003_sig000001b3
    );
  blk00000003_blk00000155 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001ba,
      Q => blk00000003_sig000001b2
    );
  blk00000003_blk00000154 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001b9,
      Q => blk00000003_sig000001b1
    );
  blk00000003_blk00000153 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001b8,
      Q => blk00000003_sig000001b0
    );
  blk00000003_blk00000152 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001b7,
      Q => blk00000003_sig000001af
    );
  blk00000003_blk00000151 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001b6,
      Q => blk00000003_sig000001ae
    );
  blk00000003_blk00000150 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001b5,
      Q => blk00000003_sig000001ad
    );
  blk00000003_blk0000014f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001b4,
      Q => blk00000003_sig000001ac
    );
  blk00000003_blk0000014e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001b3,
      Q => blk00000003_sig000001ab
    );
  blk00000003_blk0000014d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001b2,
      Q => blk00000003_sig000001aa
    );
  blk00000003_blk0000014c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001b1,
      Q => blk00000003_sig000001a9
    );
  blk00000003_blk0000014b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001b0,
      Q => blk00000003_sig000001a8
    );
  blk00000003_blk0000014a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001af,
      Q => blk00000003_sig000001a7
    );
  blk00000003_blk00000149 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001ae,
      Q => blk00000003_sig000001a6
    );
  blk00000003_blk00000148 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001ad,
      Q => blk00000003_sig000001a5
    );
  blk00000003_blk00000147 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001ac,
      Q => blk00000003_sig000001a4
    );
  blk00000003_blk00000146 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001ab,
      Q => blk00000003_sig000001a3
    );
  blk00000003_blk00000145 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001aa,
      Q => blk00000003_sig000001a2
    );
  blk00000003_blk00000144 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001a9,
      Q => blk00000003_sig000001a1
    );
  blk00000003_blk00000143 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001a8,
      Q => blk00000003_sig000001a0
    );
  blk00000003_blk00000142 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001a7,
      Q => blk00000003_sig0000019f
    );
  blk00000003_blk00000141 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001a6,
      Q => blk00000003_sig0000019e
    );
  blk00000003_blk00000140 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001a5,
      Q => blk00000003_sig0000019d
    );
  blk00000003_blk0000013f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001a4,
      Q => blk00000003_sig0000019c
    );
  blk00000003_blk0000013e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001a3,
      Q => blk00000003_sig0000019b
    );
  blk00000003_blk0000013d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001a2,
      Q => blk00000003_sig0000019a
    );
  blk00000003_blk0000013c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001a1,
      Q => blk00000003_sig00000199
    );
  blk00000003_blk0000013b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001a0,
      Q => blk00000003_sig00000198
    );
  blk00000003_blk0000013a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000019f,
      Q => blk00000003_sig00000197
    );
  blk00000003_blk00000139 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000019e,
      Q => blk00000003_sig00000196
    );
  blk00000003_blk00000138 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000019d,
      Q => blk00000003_sig00000195
    );
  blk00000003_blk00000137 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000019c,
      Q => blk00000003_sig00000194
    );
  blk00000003_blk00000136 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000019b,
      Q => blk00000003_sig00000193
    );
  blk00000003_blk00000135 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000019a,
      Q => blk00000003_sig00000192
    );
  blk00000003_blk00000134 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000199,
      Q => blk00000003_sig00000191
    );
  blk00000003_blk00000133 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000198,
      Q => blk00000003_sig00000190
    );
  blk00000003_blk00000132 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000197,
      Q => blk00000003_sig0000018f
    );
  blk00000003_blk00000131 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000196,
      Q => blk00000003_sig0000018e
    );
  blk00000003_blk00000130 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000195,
      Q => blk00000003_sig0000018d
    );
  blk00000003_blk0000012f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000194,
      Q => blk00000003_sig0000018c
    );
  blk00000003_blk0000012e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000193,
      Q => blk00000003_sig0000018b
    );
  blk00000003_blk0000012d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000192,
      Q => blk00000003_sig0000018a
    );
  blk00000003_blk0000012c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000191,
      Q => blk00000003_sig00000189
    );
  blk00000003_blk0000012b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000190,
      Q => blk00000003_sig00000188
    );
  blk00000003_blk0000012a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000018f,
      Q => blk00000003_sig00000187
    );
  blk00000003_blk00000129 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000018e,
      Q => blk00000003_sig00000186
    );
  blk00000003_blk00000128 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000018d,
      Q => blk00000003_sig00000185
    );
  blk00000003_blk00000127 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000018c,
      Q => blk00000003_sig00000184
    );
  blk00000003_blk00000126 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000018b,
      Q => blk00000003_sig00000183
    );
  blk00000003_blk00000125 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000018a,
      Q => blk00000003_sig00000182
    );
  blk00000003_blk00000124 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000189,
      Q => blk00000003_sig00000181
    );
  blk00000003_blk00000123 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000188,
      Q => blk00000003_sig00000180
    );
  blk00000003_blk00000122 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000187,
      Q => blk00000003_sig0000017f
    );
  blk00000003_blk00000121 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000186,
      Q => blk00000003_sig0000017e
    );
  blk00000003_blk00000120 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000185,
      Q => blk00000003_sig0000017d
    );
  blk00000003_blk0000011f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000184,
      Q => blk00000003_sig0000017c
    );
  blk00000003_blk0000011e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000183,
      Q => blk00000003_sig0000017b
    );
  blk00000003_blk0000011d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000182,
      Q => blk00000003_sig0000017a
    );
  blk00000003_blk0000011c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000181,
      Q => blk00000003_sig00000179
    );
  blk00000003_blk0000011b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000180,
      Q => blk00000003_sig00000178
    );
  blk00000003_blk0000011a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000017f,
      Q => blk00000003_sig00000177
    );
  blk00000003_blk00000119 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000017e,
      Q => blk00000003_sig00000176
    );
  blk00000003_blk00000118 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000017d,
      Q => blk00000003_sig00000175
    );
  blk00000003_blk00000117 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000017c,
      Q => blk00000003_sig00000174
    );
  blk00000003_blk00000116 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000017b,
      Q => blk00000003_sig00000173
    );
  blk00000003_blk00000115 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000017a,
      Q => blk00000003_sig00000172
    );
  blk00000003_blk00000114 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000179,
      Q => blk00000003_sig00000171
    );
  blk00000003_blk00000113 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000178,
      Q => blk00000003_sig00000170
    );
  blk00000003_blk00000112 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000177,
      Q => blk00000003_sig0000016f
    );
  blk00000003_blk00000111 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000176,
      Q => blk00000003_sig0000016e
    );
  blk00000003_blk00000110 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000175,
      Q => blk00000003_sig0000016d
    );
  blk00000003_blk0000010f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000174,
      Q => blk00000003_sig0000016c
    );
  blk00000003_blk0000010e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000173,
      Q => blk00000003_sig0000016b
    );
  blk00000003_blk0000010d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000172,
      Q => blk00000003_sig0000016a
    );
  blk00000003_blk0000010c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000171,
      Q => blk00000003_sig00000169
    );
  blk00000003_blk0000010b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000170,
      Q => blk00000003_sig00000168
    );
  blk00000003_blk0000010a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000016f,
      Q => blk00000003_sig00000167
    );
  blk00000003_blk00000109 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000016e,
      Q => blk00000003_sig00000166
    );
  blk00000003_blk00000108 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000016d,
      Q => blk00000003_sig00000165
    );
  blk00000003_blk00000107 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000016c,
      Q => blk00000003_sig00000164
    );
  blk00000003_blk00000106 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000016b,
      Q => blk00000003_sig00000163
    );
  blk00000003_blk00000105 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000016a,
      Q => blk00000003_sig00000162
    );
  blk00000003_blk00000104 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000169,
      Q => blk00000003_sig00000161
    );
  blk00000003_blk00000103 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000168,
      Q => blk00000003_sig00000160
    );
  blk00000003_blk00000102 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000167,
      Q => blk00000003_sig0000015f
    );
  blk00000003_blk00000101 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000166,
      Q => blk00000003_sig0000015e
    );
  blk00000003_blk00000100 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000165,
      Q => blk00000003_sig0000015d
    );
  blk00000003_blk000000ff : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000164,
      Q => blk00000003_sig0000015c
    );
  blk00000003_blk000000fe : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000163,
      Q => blk00000003_sig0000015b
    );
  blk00000003_blk000000fd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000162,
      Q => blk00000003_sig0000015a
    );
  blk00000003_blk000000fc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000161,
      Q => blk00000003_sig00000159
    );
  blk00000003_blk000000fb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000160,
      Q => blk00000003_sig00000158
    );
  blk00000003_blk000000fa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000015f,
      Q => blk00000003_sig00000157
    );
  blk00000003_blk000000f9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000015e,
      Q => blk00000003_sig00000156
    );
  blk00000003_blk000000f8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000015d,
      Q => blk00000003_sig00000155
    );
  blk00000003_blk000000f7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000015c,
      Q => blk00000003_sig00000154
    );
  blk00000003_blk000000f6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000015b,
      Q => blk00000003_sig00000153
    );
  blk00000003_blk000000f5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000015a,
      Q => blk00000003_sig00000152
    );
  blk00000003_blk000000f4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000159,
      Q => blk00000003_sig00000151
    );
  blk00000003_blk000000f3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000158,
      Q => blk00000003_sig00000150
    );
  blk00000003_blk000000f2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000157,
      Q => blk00000003_sig0000014f
    );
  blk00000003_blk000000f1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000156,
      Q => blk00000003_sig0000014e
    );
  blk00000003_blk000000f0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000155,
      Q => blk00000003_sig0000014d
    );
  blk00000003_blk000000ef : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000154,
      Q => blk00000003_sig0000014c
    );
  blk00000003_blk000000ee : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000153,
      Q => blk00000003_sig0000014b
    );
  blk00000003_blk000000ed : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000152,
      Q => blk00000003_sig0000014a
    );
  blk00000003_blk000000ec : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000151,
      Q => blk00000003_sig00000149
    );
  blk00000003_blk000000eb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000150,
      Q => blk00000003_sig00000148
    );
  blk00000003_blk000000ea : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000014f,
      Q => blk00000003_sig00000147
    );
  blk00000003_blk000000e9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000014e,
      Q => blk00000003_sig00000146
    );
  blk00000003_blk000000e8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000014d,
      Q => blk00000003_sig00000145
    );
  blk00000003_blk000000e7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000014c,
      Q => blk00000003_sig00000144
    );
  blk00000003_blk000000e6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000014b,
      Q => blk00000003_sig00000143
    );
  blk00000003_blk000000e5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000014a,
      Q => blk00000003_sig00000142
    );
  blk00000003_blk000000e4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000149,
      Q => blk00000003_sig00000141
    );
  blk00000003_blk000000e3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000148,
      Q => blk00000003_sig00000140
    );
  blk00000003_blk000000e2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000147,
      Q => blk00000003_sig0000013f
    );
  blk00000003_blk000000e1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000146,
      Q => blk00000003_sig0000013e
    );
  blk00000003_blk000000e0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000145,
      Q => blk00000003_sig0000013d
    );
  blk00000003_blk000000df : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000144,
      Q => blk00000003_sig0000013c
    );
  blk00000003_blk000000de : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000143,
      Q => blk00000003_sig0000013b
    );
  blk00000003_blk000000dd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000142,
      Q => blk00000003_sig0000013a
    );
  blk00000003_blk000000dc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000141,
      Q => blk00000003_sig00000139
    );
  blk00000003_blk000000db : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000140,
      Q => blk00000003_sig00000138
    );
  blk00000003_blk000000da : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000013f,
      Q => blk00000003_sig00000137
    );
  blk00000003_blk000000d9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000013e,
      Q => blk00000003_sig00000136
    );
  blk00000003_blk000000d8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000013d,
      Q => blk00000003_sig00000135
    );
  blk00000003_blk000000d7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000013c,
      Q => blk00000003_sig00000134
    );
  blk00000003_blk000000d6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000013b,
      Q => blk00000003_sig00000133
    );
  blk00000003_blk000000d5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000013a,
      Q => blk00000003_sig00000132
    );
  blk00000003_blk000000d4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000139,
      Q => blk00000003_sig00000131
    );
  blk00000003_blk000000d3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000138,
      Q => blk00000003_sig00000130
    );
  blk00000003_blk000000d2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000137,
      Q => blk00000003_sig0000012f
    );
  blk00000003_blk000000d1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000136,
      Q => blk00000003_sig0000012e
    );
  blk00000003_blk000000d0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000135,
      Q => blk00000003_sig0000012d
    );
  blk00000003_blk000000cf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000134,
      Q => blk00000003_sig0000012c
    );
  blk00000003_blk000000ce : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000133,
      Q => blk00000003_sig0000012b
    );
  blk00000003_blk000000cd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000132,
      Q => blk00000003_sig0000012a
    );
  blk00000003_blk000000cc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000131,
      Q => blk00000003_sig00000129
    );
  blk00000003_blk000000cb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000130,
      Q => blk00000003_sig00000128
    );
  blk00000003_blk000000ca : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000012f,
      Q => blk00000003_sig00000127
    );
  blk00000003_blk000000c9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000012e,
      Q => blk00000003_sig00000126
    );
  blk00000003_blk000000c8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000012d,
      Q => blk00000003_sig00000125
    );
  blk00000003_blk000000c7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000012c,
      Q => blk00000003_sig00000124
    );
  blk00000003_blk000000c6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000012b,
      Q => blk00000003_sig00000123
    );
  blk00000003_blk000000c5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000012a,
      Q => blk00000003_sig00000122
    );
  blk00000003_blk000000c4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000129,
      Q => blk00000003_sig00000121
    );
  blk00000003_blk000000c3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000128,
      Q => blk00000003_sig00000120
    );
  blk00000003_blk000000c2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000127,
      Q => blk00000003_sig0000011f
    );
  blk00000003_blk000000c1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000126,
      Q => blk00000003_sig0000011e
    );
  blk00000003_blk000000c0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000125,
      Q => blk00000003_sig0000011d
    );
  blk00000003_blk000000bf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000124,
      Q => blk00000003_sig0000011c
    );
  blk00000003_blk000000be : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000123,
      Q => blk00000003_sig0000011b
    );
  blk00000003_blk000000bd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000122,
      Q => blk00000003_sig0000011a
    );
  blk00000003_blk000000bc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000121,
      Q => blk00000003_sig00000119
    );
  blk00000003_blk000000bb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000120,
      Q => blk00000003_sig00000118
    );
  blk00000003_blk000000ba : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000011f,
      Q => blk00000003_sig00000117
    );
  blk00000003_blk000000b9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000011e,
      Q => blk00000003_sig00000116
    );
  blk00000003_blk000000b8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000011d,
      Q => blk00000003_sig00000115
    );
  blk00000003_blk000000b7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000011c,
      Q => blk00000003_sig00000114
    );
  blk00000003_blk000000b6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000011b,
      Q => blk00000003_sig00000113
    );
  blk00000003_blk000000b5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000011a,
      Q => blk00000003_sig00000112
    );
  blk00000003_blk000000b4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000119,
      Q => blk00000003_sig00000111
    );
  blk00000003_blk000000b3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000118,
      Q => blk00000003_sig00000110
    );
  blk00000003_blk000000b2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000117,
      Q => blk00000003_sig0000010f
    );
  blk00000003_blk000000b1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000116,
      Q => blk00000003_sig0000010e
    );
  blk00000003_blk000000b0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000115,
      Q => blk00000003_sig0000010d
    );
  blk00000003_blk000000af : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000114,
      Q => blk00000003_sig0000010c
    );
  blk00000003_blk000000ae : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000113,
      Q => blk00000003_sig0000010b
    );
  blk00000003_blk000000ad : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000112,
      Q => blk00000003_sig0000010a
    );
  blk00000003_blk000000ac : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000111,
      Q => blk00000003_sig00000109
    );
  blk00000003_blk000000ab : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000110,
      Q => blk00000003_sig00000108
    );
  blk00000003_blk000000aa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000010f,
      Q => blk00000003_sig00000107
    );
  blk00000003_blk000000a9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000010e,
      Q => blk00000003_sig00000106
    );
  blk00000003_blk000000a8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000010d,
      Q => blk00000003_sig00000105
    );
  blk00000003_blk000000a7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000010c,
      Q => blk00000003_sig00000104
    );
  blk00000003_blk000000a6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000010b,
      Q => blk00000003_sig00000103
    );
  blk00000003_blk000000a5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000010a,
      Q => blk00000003_sig00000102
    );
  blk00000003_blk000000a4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000109,
      Q => blk00000003_sig00000101
    );
  blk00000003_blk000000a3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000108,
      Q => blk00000003_sig00000100
    );
  blk00000003_blk000000a2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000107,
      Q => blk00000003_sig000000ff
    );
  blk00000003_blk000000a1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000106,
      Q => blk00000003_sig000000fe
    );
  blk00000003_blk000000a0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000105,
      Q => blk00000003_sig000000fd
    );
  blk00000003_blk0000009f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000104,
      Q => blk00000003_sig000000fc
    );
  blk00000003_blk0000009e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000103,
      Q => blk00000003_sig000000fb
    );
  blk00000003_blk0000009d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000102,
      Q => blk00000003_sig000000fa
    );
  blk00000003_blk0000009c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000101,
      Q => blk00000003_sig000000f9
    );
  blk00000003_blk0000009b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000100,
      Q => blk00000003_sig000000f8
    );
  blk00000003_blk0000009a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ff,
      Q => blk00000003_sig000000f7
    );
  blk00000003_blk00000099 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000fe,
      Q => blk00000003_sig000000f6
    );
  blk00000003_blk00000098 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000fd,
      Q => blk00000003_sig000000f5
    );
  blk00000003_blk00000097 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000fc,
      Q => blk00000003_sig000000f4
    );
  blk00000003_blk00000096 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000fb,
      Q => blk00000003_sig000000f3
    );
  blk00000003_blk00000095 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000fa,
      Q => blk00000003_sig000000f2
    );
  blk00000003_blk00000094 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f9,
      Q => blk00000003_sig000000f1
    );
  blk00000003_blk00000093 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f8,
      Q => blk00000003_sig000000f0
    );
  blk00000003_blk00000092 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f7,
      Q => blk00000003_sig000000ef
    );
  blk00000003_blk00000091 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f6,
      Q => blk00000003_sig000000ee
    );
  blk00000003_blk00000090 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f5,
      Q => blk00000003_sig000000ed
    );
  blk00000003_blk0000008f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f4,
      Q => blk00000003_sig000000ec
    );
  blk00000003_blk0000008e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f3,
      Q => blk00000003_sig000000eb
    );
  blk00000003_blk0000008d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f2,
      Q => blk00000003_sig000000e9
    );
  blk00000003_blk0000008c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f1,
      Q => blk00000003_sig000000e7
    );
  blk00000003_blk0000008b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f0,
      Q => blk00000003_sig000000e5
    );
  blk00000003_blk0000008a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ef,
      Q => blk00000003_sig000000e3
    );
  blk00000003_blk00000089 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ee,
      Q => blk00000003_sig000000e1
    );
  blk00000003_blk00000088 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ed,
      Q => blk00000003_sig000000df
    );
  blk00000003_blk00000087 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ec,
      Q => blk00000003_sig000000dd
    );
  blk00000003_blk00000086 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000eb,
      Q => blk00000003_sig000000db
    );
  blk00000003_blk00000085 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e9,
      Q => blk00000003_sig000000ea
    );
  blk00000003_blk00000084 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e7,
      Q => blk00000003_sig000000e8
    );
  blk00000003_blk00000083 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e5,
      Q => blk00000003_sig000000e6
    );
  blk00000003_blk00000082 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e3,
      Q => blk00000003_sig000000e4
    );
  blk00000003_blk00000081 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e1,
      Q => blk00000003_sig000000e2
    );
  blk00000003_blk00000080 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000df,
      Q => blk00000003_sig000000e0
    );
  blk00000003_blk0000007f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000dd,
      Q => blk00000003_sig000000de
    );
  blk00000003_blk0000007e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000db,
      Q => blk00000003_sig000000dc
    );
  blk00000003_blk0000007d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(0),
      Q => blk00000003_sig000000da
    );
  blk00000003_blk0000007c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(1),
      Q => blk00000003_sig000000d9
    );
  blk00000003_blk0000007b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(2),
      Q => blk00000003_sig000000d8
    );
  blk00000003_blk0000007a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(3),
      Q => blk00000003_sig000000d7
    );
  blk00000003_blk00000079 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(4),
      Q => blk00000003_sig000000d6
    );
  blk00000003_blk00000078 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(5),
      Q => blk00000003_sig000000d5
    );
  blk00000003_blk00000077 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(6),
      Q => blk00000003_sig000000d4
    );
  blk00000003_blk00000076 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(7),
      Q => blk00000003_sig000000d3
    );
  blk00000003_blk00000075 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(8),
      Q => blk00000003_sig000000d2
    );
  blk00000003_blk00000074 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(9),
      Q => blk00000003_sig000000d1
    );
  blk00000003_blk00000073 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(10),
      Q => blk00000003_sig000000d0
    );
  blk00000003_blk00000072 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(11),
      Q => blk00000003_sig000000cf
    );
  blk00000003_blk00000071 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(12),
      Q => blk00000003_sig000000ce
    );
  blk00000003_blk00000070 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(13),
      Q => blk00000003_sig000000cd
    );
  blk00000003_blk0000006f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(14),
      Q => blk00000003_sig000000cc
    );
  blk00000003_blk0000006e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(15),
      Q => blk00000003_sig000000cb
    );
  blk00000003_blk0000006d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(16),
      Q => blk00000003_sig000000ca
    );
  blk00000003_blk0000006c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(17),
      Q => blk00000003_sig000000c9
    );
  blk00000003_blk0000006b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(18),
      Q => blk00000003_sig000000c8
    );
  blk00000003_blk0000006a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(19),
      Q => blk00000003_sig000000c7
    );
  blk00000003_blk00000069 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(20),
      Q => blk00000003_sig000000c6
    );
  blk00000003_blk00000068 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(21),
      Q => blk00000003_sig000000c5
    );
  blk00000003_blk00000067 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(22),
      Q => blk00000003_sig000000c4
    );
  blk00000003_blk00000066 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(23),
      Q => blk00000003_sig000000c3
    );
  blk00000003_blk00000065 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(24),
      Q => blk00000003_sig000000c2
    );
  blk00000003_blk00000064 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(25),
      Q => blk00000003_sig000000c1
    );
  blk00000003_blk00000063 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(26),
      Q => blk00000003_sig000000c0
    );
  blk00000003_blk00000062 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(27),
      Q => blk00000003_sig000000bf
    );
  blk00000003_blk00000061 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(28),
      Q => blk00000003_sig000000be
    );
  blk00000003_blk00000060 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(29),
      Q => blk00000003_sig000000bd
    );
  blk00000003_blk0000005f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(30),
      Q => blk00000003_sig000000bc
    );
  blk00000003_blk0000005e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(31),
      Q => blk00000003_sig000000bb
    );
  blk00000003_blk0000005d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ba,
      Q => quotient(0)
    );
  blk00000003_blk0000005c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b9,
      Q => quotient(1)
    );
  blk00000003_blk0000005b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b8,
      Q => quotient(2)
    );
  blk00000003_blk0000005a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b7,
      Q => quotient(3)
    );
  blk00000003_blk00000059 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b6,
      Q => quotient(4)
    );
  blk00000003_blk00000058 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b5,
      Q => quotient(5)
    );
  blk00000003_blk00000057 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b4,
      Q => quotient(6)
    );
  blk00000003_blk00000056 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b3,
      Q => quotient(7)
    );
  blk00000003_blk00000055 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b2,
      Q => quotient(8)
    );
  blk00000003_blk00000054 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b1,
      Q => quotient(9)
    );
  blk00000003_blk00000053 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b0,
      Q => quotient(10)
    );
  blk00000003_blk00000052 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000af,
      Q => quotient(11)
    );
  blk00000003_blk00000051 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ae,
      Q => quotient(12)
    );
  blk00000003_blk00000050 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ad,
      Q => quotient(13)
    );
  blk00000003_blk0000004f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ac,
      Q => quotient(14)
    );
  blk00000003_blk0000004e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ab,
      Q => quotient(15)
    );
  blk00000003_blk0000004d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000aa,
      Q => quotient(16)
    );
  blk00000003_blk0000004c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a9,
      Q => quotient(17)
    );
  blk00000003_blk0000004b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a8,
      Q => quotient(18)
    );
  blk00000003_blk0000004a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a7,
      Q => quotient(19)
    );
  blk00000003_blk00000049 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a6,
      Q => quotient(20)
    );
  blk00000003_blk00000048 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a5,
      Q => quotient(21)
    );
  blk00000003_blk00000047 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a4,
      Q => quotient(22)
    );
  blk00000003_blk00000046 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a3,
      Q => quotient(23)
    );
  blk00000003_blk00000045 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a2,
      Q => quotient(24)
    );
  blk00000003_blk00000044 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a1,
      Q => quotient(25)
    );
  blk00000003_blk00000043 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a0,
      Q => quotient(26)
    );
  blk00000003_blk00000042 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000009f,
      Q => quotient(27)
    );
  blk00000003_blk00000041 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000009e,
      Q => quotient(28)
    );
  blk00000003_blk00000040 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000009d,
      Q => quotient(29)
    );
  blk00000003_blk0000003f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000009c,
      Q => quotient(30)
    );
  blk00000003_blk0000003e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000009b,
      Q => quotient(31)
    );
  blk00000003_blk0000003d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000056,
      Q => blk00000003_sig0000009a
    );
  blk00000003_blk0000003c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000099,
      Q => blk00000003_sig00000098
    );
  blk00000003_blk0000003b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000098,
      Q => blk00000003_sig00000096
    );
  blk00000003_blk0000003a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000097,
      Q => blk00000003_sig00000095
    );
  blk00000003_blk00000039 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000096,
      Q => blk00000003_sig00000093
    );
  blk00000003_blk00000038 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000095,
      Q => blk00000003_sig00000092
    );
  blk00000003_blk00000037 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000094,
      Q => blk00000003_sig00000091
    );
  blk00000003_blk00000036 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000093,
      Q => blk00000003_sig0000008f
    );
  blk00000003_blk00000035 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000092,
      Q => blk00000003_sig0000008e
    );
  blk00000003_blk00000034 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000091,
      Q => blk00000003_sig0000008d
    );
  blk00000003_blk00000033 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000090,
      Q => blk00000003_sig0000008c
    );
  blk00000003_blk00000032 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000008f,
      Q => blk00000003_sig0000008a
    );
  blk00000003_blk00000031 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000008e,
      Q => blk00000003_sig00000089
    );
  blk00000003_blk00000030 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000008d,
      Q => blk00000003_sig00000088
    );
  blk00000003_blk0000002f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000008c,
      Q => blk00000003_sig00000087
    );
  blk00000003_blk0000002e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000008b,
      Q => blk00000003_sig00000086
    );
  blk00000003_blk0000002d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000008a,
      Q => blk00000003_sig00000083
    );
  blk00000003_blk0000002c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000089,
      Q => blk00000003_sig00000081
    );
  blk00000003_blk0000002b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000088,
      Q => blk00000003_sig0000007f
    );
  blk00000003_blk0000002a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000087,
      Q => blk00000003_sig0000007d
    );
  blk00000003_blk00000029 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000086,
      Q => blk00000003_sig0000007b
    );
  blk00000003_blk00000028 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000085,
      Q => blk00000003_sig00000079
    );
  blk00000003_blk00000027 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000083,
      Q => blk00000003_sig00000084
    );
  blk00000003_blk00000026 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000081,
      Q => blk00000003_sig00000082
    );
  blk00000003_blk00000025 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007f,
      Q => blk00000003_sig00000080
    );
  blk00000003_blk00000024 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007d,
      Q => blk00000003_sig0000007e
    );
  blk00000003_blk00000023 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007b,
      Q => blk00000003_sig0000007c
    );
  blk00000003_blk00000022 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000079,
      Q => blk00000003_sig0000007a
    );
  blk00000003_blk00000021 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000077,
      Q => blk00000003_sig00000078
    );
  blk00000003_blk00000020 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000075,
      Q => blk00000003_sig00000076
    );
  blk00000003_blk0000001f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000074,
      Q => blk00000003_sig0000006d
    );
  blk00000003_blk0000001e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000073,
      Q => blk00000003_sig0000006c
    );
  blk00000003_blk0000001d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000072,
      Q => blk00000003_sig0000006b
    );
  blk00000003_blk0000001c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000071,
      Q => blk00000003_sig0000006a
    );
  blk00000003_blk0000001b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000070,
      Q => blk00000003_sig00000069
    );
  blk00000003_blk0000001a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006f,
      Q => blk00000003_sig00000068
    );
  blk00000003_blk00000019 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006d,
      Q => blk00000003_sig0000006e
    );
  blk00000003_blk00000018 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006c,
      Q => blk00000003_sig00000066
    );
  blk00000003_blk00000017 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006b,
      Q => blk00000003_sig00000065
    );
  blk00000003_blk00000016 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006a,
      Q => blk00000003_sig00000064
    );
  blk00000003_blk00000015 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000069,
      Q => blk00000003_sig00000063
    );
  blk00000003_blk00000014 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000068,
      Q => blk00000003_sig00000062
    );
  blk00000003_blk00000013 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000066,
      Q => blk00000003_sig00000067
    );
  blk00000003_blk00000012 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000065,
      Q => blk00000003_sig00000060
    );
  blk00000003_blk00000011 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000064,
      Q => blk00000003_sig0000005f
    );
  blk00000003_blk00000010 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000063,
      Q => blk00000003_sig0000005e
    );
  blk00000003_blk0000000f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000062,
      Q => blk00000003_sig0000005d
    );
  blk00000003_blk0000000e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000060,
      Q => blk00000003_sig00000061
    );
  blk00000003_blk0000000d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000005f,
      Q => blk00000003_sig0000005b
    );
  blk00000003_blk0000000c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000005e,
      Q => blk00000003_sig0000005a
    );
  blk00000003_blk0000000b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000005d,
      Q => blk00000003_sig00000059
    );
  blk00000003_blk0000000a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000005b,
      Q => blk00000003_sig0000005c
    );
  blk00000003_blk00000009 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000005a,
      Q => blk00000003_sig00000057
    );
  blk00000003_blk00000008 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000059,
      Q => blk00000003_sig00000055
    );
  blk00000003_blk00000007 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000057,
      Q => blk00000003_sig00000058
    );
  blk00000003_blk00000006 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000055,
      Q => blk00000003_sig00000056
    );
  blk00000003_blk00000005 : VCC
    port map (
      P => NlwRenamedSig_OI_rfd
    );
  blk00000003_blk00000004 : GND
    port map (
      G => blk00000003_sig00000053
    );

end STRUCTURE;

-- synthesis translate_on
--------------------------------------------------------------------------------
-- Copyright (c) 1995-2011 Xilinx, Inc.  All rights reserved.
--------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /    Vendor: Xilinx
-- \   \   \/     Version: O.61xd
--  \   \         Application: netgen
--  /   /         Filename: dv_gn_v3_0_90662698f61d80cb.vhd
-- /___/   /\     Timestamp: Mon Jul 23 19:56:37 2012
-- \   \  /  \ 
--  \___\/\___\
--             
-- Command	: -intstyle ise -w -sim -ofmt vhdl ./tmp/_cg/dv_gn_v3_0_90662698f61d80cb.ngc ./tmp/_cg/dv_gn_v3_0_90662698f61d80cb.vhd 
-- Device	: 6vcx75tff484-2
-- Input file	: ./tmp/_cg/dv_gn_v3_0_90662698f61d80cb.ngc
-- Output file	: ./tmp/_cg/dv_gn_v3_0_90662698f61d80cb.vhd
-- # of Entities	: 1
-- Design Name	: dv_gn_v3_0_90662698f61d80cb
-- Xilinx	: c:\xilinx\13.2\ise_ds\ise\
--             
-- Purpose:    
--     This VHDL netlist is a verification model and uses simulation 
--     primitives which may not represent the true implementation of the 
--     device, however the netlist is functionally correct and should not 
--     be modified. This file cannot be synthesized and should only be used 
--     with supported simulation tools.
--             
-- Reference:  
--     Command Line Tools User Guide, Chapter 23
--     Synthesis and Simulation Design Guide, Chapter 6
--             
--------------------------------------------------------------------------------


-- synthesis translate_off
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;
use UNISIM.VPKG.ALL;

entity dv_gn_v3_0_90662698f61d80cb is
  port (
    ce : in STD_LOGIC := 'X'; 
    rfd : out STD_LOGIC; 
    clk : in STD_LOGIC := 'X'; 
    dividend : in STD_LOGIC_VECTOR ( 31 downto 0 ); 
    quotient : out STD_LOGIC_VECTOR ( 31 downto 0 ); 
    divisor : in STD_LOGIC_VECTOR ( 5 downto 0 ); 
    fractional : out STD_LOGIC_VECTOR ( 5 downto 0 ) 
  );
end dv_gn_v3_0_90662698f61d80cb;

architecture STRUCTURE of dv_gn_v3_0_90662698f61d80cb is
  signal NlwRenamedSig_OI_rfd : STD_LOGIC; 
  signal blk00000003_sig00000910 : STD_LOGIC; 
  signal blk00000003_sig0000090f : STD_LOGIC; 
  signal blk00000003_sig0000090e : STD_LOGIC; 
  signal blk00000003_sig0000090d : STD_LOGIC; 
  signal blk00000003_sig0000090c : STD_LOGIC; 
  signal blk00000003_sig0000090b : STD_LOGIC; 
  signal blk00000003_sig0000090a : STD_LOGIC; 
  signal blk00000003_sig00000909 : STD_LOGIC; 
  signal blk00000003_sig00000908 : STD_LOGIC; 
  signal blk00000003_sig00000907 : STD_LOGIC; 
  signal blk00000003_sig00000906 : STD_LOGIC; 
  signal blk00000003_sig00000905 : STD_LOGIC; 
  signal blk00000003_sig00000904 : STD_LOGIC; 
  signal blk00000003_sig00000903 : STD_LOGIC; 
  signal blk00000003_sig00000902 : STD_LOGIC; 
  signal blk00000003_sig00000901 : STD_LOGIC; 
  signal blk00000003_sig00000900 : STD_LOGIC; 
  signal blk00000003_sig000008ff : STD_LOGIC; 
  signal blk00000003_sig000008fe : STD_LOGIC; 
  signal blk00000003_sig000008fd : STD_LOGIC; 
  signal blk00000003_sig000008fc : STD_LOGIC; 
  signal blk00000003_sig000008fb : STD_LOGIC; 
  signal blk00000003_sig000008fa : STD_LOGIC; 
  signal blk00000003_sig000008f9 : STD_LOGIC; 
  signal blk00000003_sig000008f8 : STD_LOGIC; 
  signal blk00000003_sig000008f7 : STD_LOGIC; 
  signal blk00000003_sig000008f6 : STD_LOGIC; 
  signal blk00000003_sig000008f5 : STD_LOGIC; 
  signal blk00000003_sig000008f4 : STD_LOGIC; 
  signal blk00000003_sig000008f3 : STD_LOGIC; 
  signal blk00000003_sig000008f2 : STD_LOGIC; 
  signal blk00000003_sig000008f1 : STD_LOGIC; 
  signal blk00000003_sig000008f0 : STD_LOGIC; 
  signal blk00000003_sig000008ef : STD_LOGIC; 
  signal blk00000003_sig000008ee : STD_LOGIC; 
  signal blk00000003_sig000008ed : STD_LOGIC; 
  signal blk00000003_sig000008ec : STD_LOGIC; 
  signal blk00000003_sig000008eb : STD_LOGIC; 
  signal blk00000003_sig000008ea : STD_LOGIC; 
  signal blk00000003_sig000008e9 : STD_LOGIC; 
  signal blk00000003_sig000008e8 : STD_LOGIC; 
  signal blk00000003_sig000008e7 : STD_LOGIC; 
  signal blk00000003_sig000008e6 : STD_LOGIC; 
  signal blk00000003_sig000008e5 : STD_LOGIC; 
  signal blk00000003_sig000008e4 : STD_LOGIC; 
  signal blk00000003_sig000008e3 : STD_LOGIC; 
  signal blk00000003_sig000008e2 : STD_LOGIC; 
  signal blk00000003_sig000008e1 : STD_LOGIC; 
  signal blk00000003_sig000008e0 : STD_LOGIC; 
  signal blk00000003_sig000008df : STD_LOGIC; 
  signal blk00000003_sig000008de : STD_LOGIC; 
  signal blk00000003_sig000008dd : STD_LOGIC; 
  signal blk00000003_sig000008dc : STD_LOGIC; 
  signal blk00000003_sig000008db : STD_LOGIC; 
  signal blk00000003_sig000008da : STD_LOGIC; 
  signal blk00000003_sig000008d9 : STD_LOGIC; 
  signal blk00000003_sig000008d8 : STD_LOGIC; 
  signal blk00000003_sig000008d7 : STD_LOGIC; 
  signal blk00000003_sig000008d6 : STD_LOGIC; 
  signal blk00000003_sig000008d5 : STD_LOGIC; 
  signal blk00000003_sig000008d4 : STD_LOGIC; 
  signal blk00000003_sig000008d3 : STD_LOGIC; 
  signal blk00000003_sig000008d2 : STD_LOGIC; 
  signal blk00000003_sig000008d1 : STD_LOGIC; 
  signal blk00000003_sig000008d0 : STD_LOGIC; 
  signal blk00000003_sig000008cf : STD_LOGIC; 
  signal blk00000003_sig000008ce : STD_LOGIC; 
  signal blk00000003_sig000008cd : STD_LOGIC; 
  signal blk00000003_sig000008cc : STD_LOGIC; 
  signal blk00000003_sig000008cb : STD_LOGIC; 
  signal blk00000003_sig000008ca : STD_LOGIC; 
  signal blk00000003_sig000008c9 : STD_LOGIC; 
  signal blk00000003_sig000008c8 : STD_LOGIC; 
  signal blk00000003_sig000008c7 : STD_LOGIC; 
  signal blk00000003_sig000008c6 : STD_LOGIC; 
  signal blk00000003_sig000008c5 : STD_LOGIC; 
  signal blk00000003_sig000008c4 : STD_LOGIC; 
  signal blk00000003_sig000008c3 : STD_LOGIC; 
  signal blk00000003_sig000008c2 : STD_LOGIC; 
  signal blk00000003_sig000008c1 : STD_LOGIC; 
  signal blk00000003_sig000008c0 : STD_LOGIC; 
  signal blk00000003_sig000008bf : STD_LOGIC; 
  signal blk00000003_sig000008be : STD_LOGIC; 
  signal blk00000003_sig000008bd : STD_LOGIC; 
  signal blk00000003_sig000008bc : STD_LOGIC; 
  signal blk00000003_sig000008bb : STD_LOGIC; 
  signal blk00000003_sig000008ba : STD_LOGIC; 
  signal blk00000003_sig000008b9 : STD_LOGIC; 
  signal blk00000003_sig000008b8 : STD_LOGIC; 
  signal blk00000003_sig000008b7 : STD_LOGIC; 
  signal blk00000003_sig000008b6 : STD_LOGIC; 
  signal blk00000003_sig000008b5 : STD_LOGIC; 
  signal blk00000003_sig000008b4 : STD_LOGIC; 
  signal blk00000003_sig000008b3 : STD_LOGIC; 
  signal blk00000003_sig000008b2 : STD_LOGIC; 
  signal blk00000003_sig000008b1 : STD_LOGIC; 
  signal blk00000003_sig000008b0 : STD_LOGIC; 
  signal blk00000003_sig000008af : STD_LOGIC; 
  signal blk00000003_sig000008ae : STD_LOGIC; 
  signal blk00000003_sig000008ad : STD_LOGIC; 
  signal blk00000003_sig000008ac : STD_LOGIC; 
  signal blk00000003_sig000008ab : STD_LOGIC; 
  signal blk00000003_sig000008aa : STD_LOGIC; 
  signal blk00000003_sig000008a9 : STD_LOGIC; 
  signal blk00000003_sig000008a8 : STD_LOGIC; 
  signal blk00000003_sig000008a7 : STD_LOGIC; 
  signal blk00000003_sig000008a6 : STD_LOGIC; 
  signal blk00000003_sig000008a5 : STD_LOGIC; 
  signal blk00000003_sig000008a4 : STD_LOGIC; 
  signal blk00000003_sig000008a3 : STD_LOGIC; 
  signal blk00000003_sig000008a2 : STD_LOGIC; 
  signal blk00000003_sig000008a1 : STD_LOGIC; 
  signal blk00000003_sig000008a0 : STD_LOGIC; 
  signal blk00000003_sig0000089f : STD_LOGIC; 
  signal blk00000003_sig0000089e : STD_LOGIC; 
  signal blk00000003_sig0000089d : STD_LOGIC; 
  signal blk00000003_sig0000089c : STD_LOGIC; 
  signal blk00000003_sig0000089b : STD_LOGIC; 
  signal blk00000003_sig0000089a : STD_LOGIC; 
  signal blk00000003_sig00000899 : STD_LOGIC; 
  signal blk00000003_sig00000898 : STD_LOGIC; 
  signal blk00000003_sig00000897 : STD_LOGIC; 
  signal blk00000003_sig00000896 : STD_LOGIC; 
  signal blk00000003_sig00000895 : STD_LOGIC; 
  signal blk00000003_sig00000894 : STD_LOGIC; 
  signal blk00000003_sig00000893 : STD_LOGIC; 
  signal blk00000003_sig00000892 : STD_LOGIC; 
  signal blk00000003_sig00000891 : STD_LOGIC; 
  signal blk00000003_sig00000890 : STD_LOGIC; 
  signal blk00000003_sig0000088f : STD_LOGIC; 
  signal blk00000003_sig0000088e : STD_LOGIC; 
  signal blk00000003_sig0000088d : STD_LOGIC; 
  signal blk00000003_sig0000088c : STD_LOGIC; 
  signal blk00000003_sig0000088b : STD_LOGIC; 
  signal blk00000003_sig0000088a : STD_LOGIC; 
  signal blk00000003_sig00000889 : STD_LOGIC; 
  signal blk00000003_sig00000888 : STD_LOGIC; 
  signal blk00000003_sig00000887 : STD_LOGIC; 
  signal blk00000003_sig00000886 : STD_LOGIC; 
  signal blk00000003_sig00000885 : STD_LOGIC; 
  signal blk00000003_sig00000884 : STD_LOGIC; 
  signal blk00000003_sig00000883 : STD_LOGIC; 
  signal blk00000003_sig00000882 : STD_LOGIC; 
  signal blk00000003_sig00000881 : STD_LOGIC; 
  signal blk00000003_sig00000880 : STD_LOGIC; 
  signal blk00000003_sig0000087f : STD_LOGIC; 
  signal blk00000003_sig0000087e : STD_LOGIC; 
  signal blk00000003_sig0000087d : STD_LOGIC; 
  signal blk00000003_sig0000087c : STD_LOGIC; 
  signal blk00000003_sig0000087b : STD_LOGIC; 
  signal blk00000003_sig0000087a : STD_LOGIC; 
  signal blk00000003_sig00000879 : STD_LOGIC; 
  signal blk00000003_sig00000878 : STD_LOGIC; 
  signal blk00000003_sig00000877 : STD_LOGIC; 
  signal blk00000003_sig00000876 : STD_LOGIC; 
  signal blk00000003_sig00000875 : STD_LOGIC; 
  signal blk00000003_sig00000874 : STD_LOGIC; 
  signal blk00000003_sig00000873 : STD_LOGIC; 
  signal blk00000003_sig00000872 : STD_LOGIC; 
  signal blk00000003_sig00000871 : STD_LOGIC; 
  signal blk00000003_sig00000870 : STD_LOGIC; 
  signal blk00000003_sig0000086f : STD_LOGIC; 
  signal blk00000003_sig0000086e : STD_LOGIC; 
  signal blk00000003_sig0000086d : STD_LOGIC; 
  signal blk00000003_sig0000086c : STD_LOGIC; 
  signal blk00000003_sig0000086b : STD_LOGIC; 
  signal blk00000003_sig0000086a : STD_LOGIC; 
  signal blk00000003_sig00000869 : STD_LOGIC; 
  signal blk00000003_sig00000868 : STD_LOGIC; 
  signal blk00000003_sig00000867 : STD_LOGIC; 
  signal blk00000003_sig00000866 : STD_LOGIC; 
  signal blk00000003_sig00000865 : STD_LOGIC; 
  signal blk00000003_sig00000864 : STD_LOGIC; 
  signal blk00000003_sig00000863 : STD_LOGIC; 
  signal blk00000003_sig00000862 : STD_LOGIC; 
  signal blk00000003_sig00000861 : STD_LOGIC; 
  signal blk00000003_sig00000860 : STD_LOGIC; 
  signal blk00000003_sig0000085f : STD_LOGIC; 
  signal blk00000003_sig0000085e : STD_LOGIC; 
  signal blk00000003_sig0000085d : STD_LOGIC; 
  signal blk00000003_sig0000085c : STD_LOGIC; 
  signal blk00000003_sig0000085b : STD_LOGIC; 
  signal blk00000003_sig0000085a : STD_LOGIC; 
  signal blk00000003_sig00000859 : STD_LOGIC; 
  signal blk00000003_sig00000858 : STD_LOGIC; 
  signal blk00000003_sig00000857 : STD_LOGIC; 
  signal blk00000003_sig00000856 : STD_LOGIC; 
  signal blk00000003_sig00000855 : STD_LOGIC; 
  signal blk00000003_sig00000854 : STD_LOGIC; 
  signal blk00000003_sig00000853 : STD_LOGIC; 
  signal blk00000003_sig00000852 : STD_LOGIC; 
  signal blk00000003_sig00000851 : STD_LOGIC; 
  signal blk00000003_sig00000850 : STD_LOGIC; 
  signal blk00000003_sig0000084f : STD_LOGIC; 
  signal blk00000003_sig0000084e : STD_LOGIC; 
  signal blk00000003_sig0000084d : STD_LOGIC; 
  signal blk00000003_sig0000084c : STD_LOGIC; 
  signal blk00000003_sig0000084b : STD_LOGIC; 
  signal blk00000003_sig0000084a : STD_LOGIC; 
  signal blk00000003_sig00000849 : STD_LOGIC; 
  signal blk00000003_sig00000848 : STD_LOGIC; 
  signal blk00000003_sig00000847 : STD_LOGIC; 
  signal blk00000003_sig00000846 : STD_LOGIC; 
  signal blk00000003_sig00000845 : STD_LOGIC; 
  signal blk00000003_sig00000844 : STD_LOGIC; 
  signal blk00000003_sig00000843 : STD_LOGIC; 
  signal blk00000003_sig00000842 : STD_LOGIC; 
  signal blk00000003_sig00000841 : STD_LOGIC; 
  signal blk00000003_sig00000840 : STD_LOGIC; 
  signal blk00000003_sig0000083f : STD_LOGIC; 
  signal blk00000003_sig0000083e : STD_LOGIC; 
  signal blk00000003_sig0000083d : STD_LOGIC; 
  signal blk00000003_sig0000083c : STD_LOGIC; 
  signal blk00000003_sig0000083b : STD_LOGIC; 
  signal blk00000003_sig0000083a : STD_LOGIC; 
  signal blk00000003_sig00000839 : STD_LOGIC; 
  signal blk00000003_sig00000838 : STD_LOGIC; 
  signal blk00000003_sig00000837 : STD_LOGIC; 
  signal blk00000003_sig00000836 : STD_LOGIC; 
  signal blk00000003_sig00000835 : STD_LOGIC; 
  signal blk00000003_sig00000834 : STD_LOGIC; 
  signal blk00000003_sig00000833 : STD_LOGIC; 
  signal blk00000003_sig00000832 : STD_LOGIC; 
  signal blk00000003_sig00000831 : STD_LOGIC; 
  signal blk00000003_sig00000830 : STD_LOGIC; 
  signal blk00000003_sig0000082f : STD_LOGIC; 
  signal blk00000003_sig0000082e : STD_LOGIC; 
  signal blk00000003_sig0000082d : STD_LOGIC; 
  signal blk00000003_sig0000082c : STD_LOGIC; 
  signal blk00000003_sig0000082b : STD_LOGIC; 
  signal blk00000003_sig0000082a : STD_LOGIC; 
  signal blk00000003_sig00000829 : STD_LOGIC; 
  signal blk00000003_sig00000828 : STD_LOGIC; 
  signal blk00000003_sig00000827 : STD_LOGIC; 
  signal blk00000003_sig00000826 : STD_LOGIC; 
  signal blk00000003_sig00000825 : STD_LOGIC; 
  signal blk00000003_sig00000824 : STD_LOGIC; 
  signal blk00000003_sig00000823 : STD_LOGIC; 
  signal blk00000003_sig00000822 : STD_LOGIC; 
  signal blk00000003_sig00000821 : STD_LOGIC; 
  signal blk00000003_sig00000820 : STD_LOGIC; 
  signal blk00000003_sig0000081f : STD_LOGIC; 
  signal blk00000003_sig0000081e : STD_LOGIC; 
  signal blk00000003_sig0000081d : STD_LOGIC; 
  signal blk00000003_sig0000081c : STD_LOGIC; 
  signal blk00000003_sig0000081b : STD_LOGIC; 
  signal blk00000003_sig0000081a : STD_LOGIC; 
  signal blk00000003_sig00000819 : STD_LOGIC; 
  signal blk00000003_sig00000818 : STD_LOGIC; 
  signal blk00000003_sig00000817 : STD_LOGIC; 
  signal blk00000003_sig00000816 : STD_LOGIC; 
  signal blk00000003_sig00000815 : STD_LOGIC; 
  signal blk00000003_sig00000814 : STD_LOGIC; 
  signal blk00000003_sig00000813 : STD_LOGIC; 
  signal blk00000003_sig00000812 : STD_LOGIC; 
  signal blk00000003_sig00000811 : STD_LOGIC; 
  signal blk00000003_sig00000810 : STD_LOGIC; 
  signal blk00000003_sig0000080f : STD_LOGIC; 
  signal blk00000003_sig0000080e : STD_LOGIC; 
  signal blk00000003_sig0000080d : STD_LOGIC; 
  signal blk00000003_sig0000080c : STD_LOGIC; 
  signal blk00000003_sig0000080b : STD_LOGIC; 
  signal blk00000003_sig0000080a : STD_LOGIC; 
  signal blk00000003_sig00000809 : STD_LOGIC; 
  signal blk00000003_sig00000808 : STD_LOGIC; 
  signal blk00000003_sig00000807 : STD_LOGIC; 
  signal blk00000003_sig00000806 : STD_LOGIC; 
  signal blk00000003_sig00000805 : STD_LOGIC; 
  signal blk00000003_sig00000804 : STD_LOGIC; 
  signal blk00000003_sig00000803 : STD_LOGIC; 
  signal blk00000003_sig00000802 : STD_LOGIC; 
  signal blk00000003_sig00000801 : STD_LOGIC; 
  signal blk00000003_sig00000800 : STD_LOGIC; 
  signal blk00000003_sig000007ff : STD_LOGIC; 
  signal blk00000003_sig000007fe : STD_LOGIC; 
  signal blk00000003_sig000007fd : STD_LOGIC; 
  signal blk00000003_sig000007fc : STD_LOGIC; 
  signal blk00000003_sig000007fb : STD_LOGIC; 
  signal blk00000003_sig000007fa : STD_LOGIC; 
  signal blk00000003_sig000007f9 : STD_LOGIC; 
  signal blk00000003_sig000007f8 : STD_LOGIC; 
  signal blk00000003_sig000007f7 : STD_LOGIC; 
  signal blk00000003_sig000007f6 : STD_LOGIC; 
  signal blk00000003_sig000007f5 : STD_LOGIC; 
  signal blk00000003_sig000007f4 : STD_LOGIC; 
  signal blk00000003_sig000007f3 : STD_LOGIC; 
  signal blk00000003_sig000007f2 : STD_LOGIC; 
  signal blk00000003_sig000007f1 : STD_LOGIC; 
  signal blk00000003_sig000007f0 : STD_LOGIC; 
  signal blk00000003_sig000007ef : STD_LOGIC; 
  signal blk00000003_sig000007ee : STD_LOGIC; 
  signal blk00000003_sig000007ed : STD_LOGIC; 
  signal blk00000003_sig000007ec : STD_LOGIC; 
  signal blk00000003_sig000007eb : STD_LOGIC; 
  signal blk00000003_sig000007ea : STD_LOGIC; 
  signal blk00000003_sig000007e9 : STD_LOGIC; 
  signal blk00000003_sig000007e8 : STD_LOGIC; 
  signal blk00000003_sig000007e7 : STD_LOGIC; 
  signal blk00000003_sig000007e6 : STD_LOGIC; 
  signal blk00000003_sig000007e5 : STD_LOGIC; 
  signal blk00000003_sig000007e4 : STD_LOGIC; 
  signal blk00000003_sig000007e3 : STD_LOGIC; 
  signal blk00000003_sig000007e2 : STD_LOGIC; 
  signal blk00000003_sig000007e1 : STD_LOGIC; 
  signal blk00000003_sig000007e0 : STD_LOGIC; 
  signal blk00000003_sig000007df : STD_LOGIC; 
  signal blk00000003_sig000007de : STD_LOGIC; 
  signal blk00000003_sig000007dd : STD_LOGIC; 
  signal blk00000003_sig000007dc : STD_LOGIC; 
  signal blk00000003_sig000007db : STD_LOGIC; 
  signal blk00000003_sig000007da : STD_LOGIC; 
  signal blk00000003_sig000007d9 : STD_LOGIC; 
  signal blk00000003_sig000007d8 : STD_LOGIC; 
  signal blk00000003_sig000007d7 : STD_LOGIC; 
  signal blk00000003_sig000007d6 : STD_LOGIC; 
  signal blk00000003_sig000007d5 : STD_LOGIC; 
  signal blk00000003_sig000007d4 : STD_LOGIC; 
  signal blk00000003_sig000007d3 : STD_LOGIC; 
  signal blk00000003_sig000007d2 : STD_LOGIC; 
  signal blk00000003_sig000007d1 : STD_LOGIC; 
  signal blk00000003_sig000007d0 : STD_LOGIC; 
  signal blk00000003_sig000007cf : STD_LOGIC; 
  signal blk00000003_sig000007ce : STD_LOGIC; 
  signal blk00000003_sig000007cd : STD_LOGIC; 
  signal blk00000003_sig000007cc : STD_LOGIC; 
  signal blk00000003_sig000007cb : STD_LOGIC; 
  signal blk00000003_sig000007ca : STD_LOGIC; 
  signal blk00000003_sig000007c9 : STD_LOGIC; 
  signal blk00000003_sig000007c8 : STD_LOGIC; 
  signal blk00000003_sig000007c7 : STD_LOGIC; 
  signal blk00000003_sig000007c6 : STD_LOGIC; 
  signal blk00000003_sig000007c5 : STD_LOGIC; 
  signal blk00000003_sig000007c4 : STD_LOGIC; 
  signal blk00000003_sig000007c3 : STD_LOGIC; 
  signal blk00000003_sig000007c2 : STD_LOGIC; 
  signal blk00000003_sig000007c1 : STD_LOGIC; 
  signal blk00000003_sig000007c0 : STD_LOGIC; 
  signal blk00000003_sig000007bf : STD_LOGIC; 
  signal blk00000003_sig000007be : STD_LOGIC; 
  signal blk00000003_sig000007bd : STD_LOGIC; 
  signal blk00000003_sig000007bc : STD_LOGIC; 
  signal blk00000003_sig000007bb : STD_LOGIC; 
  signal blk00000003_sig000007ba : STD_LOGIC; 
  signal blk00000003_sig000007b9 : STD_LOGIC; 
  signal blk00000003_sig000007b8 : STD_LOGIC; 
  signal blk00000003_sig000007b7 : STD_LOGIC; 
  signal blk00000003_sig000007b6 : STD_LOGIC; 
  signal blk00000003_sig000007b5 : STD_LOGIC; 
  signal blk00000003_sig000007b4 : STD_LOGIC; 
  signal blk00000003_sig000007b3 : STD_LOGIC; 
  signal blk00000003_sig000007b2 : STD_LOGIC; 
  signal blk00000003_sig000007b1 : STD_LOGIC; 
  signal blk00000003_sig000007b0 : STD_LOGIC; 
  signal blk00000003_sig000007af : STD_LOGIC; 
  signal blk00000003_sig000007ae : STD_LOGIC; 
  signal blk00000003_sig000007ad : STD_LOGIC; 
  signal blk00000003_sig000007ac : STD_LOGIC; 
  signal blk00000003_sig000007ab : STD_LOGIC; 
  signal blk00000003_sig000007aa : STD_LOGIC; 
  signal blk00000003_sig000007a9 : STD_LOGIC; 
  signal blk00000003_sig000007a8 : STD_LOGIC; 
  signal blk00000003_sig000007a7 : STD_LOGIC; 
  signal blk00000003_sig000007a6 : STD_LOGIC; 
  signal blk00000003_sig000007a5 : STD_LOGIC; 
  signal blk00000003_sig000007a4 : STD_LOGIC; 
  signal blk00000003_sig000007a3 : STD_LOGIC; 
  signal blk00000003_sig000007a2 : STD_LOGIC; 
  signal blk00000003_sig000007a1 : STD_LOGIC; 
  signal blk00000003_sig000007a0 : STD_LOGIC; 
  signal blk00000003_sig0000079f : STD_LOGIC; 
  signal blk00000003_sig0000079e : STD_LOGIC; 
  signal blk00000003_sig0000079d : STD_LOGIC; 
  signal blk00000003_sig0000079c : STD_LOGIC; 
  signal blk00000003_sig0000079b : STD_LOGIC; 
  signal blk00000003_sig0000079a : STD_LOGIC; 
  signal blk00000003_sig00000799 : STD_LOGIC; 
  signal blk00000003_sig00000798 : STD_LOGIC; 
  signal blk00000003_sig00000797 : STD_LOGIC; 
  signal blk00000003_sig00000796 : STD_LOGIC; 
  signal blk00000003_sig00000795 : STD_LOGIC; 
  signal blk00000003_sig00000794 : STD_LOGIC; 
  signal blk00000003_sig00000793 : STD_LOGIC; 
  signal blk00000003_sig00000792 : STD_LOGIC; 
  signal blk00000003_sig00000791 : STD_LOGIC; 
  signal blk00000003_sig00000790 : STD_LOGIC; 
  signal blk00000003_sig0000078f : STD_LOGIC; 
  signal blk00000003_sig0000078e : STD_LOGIC; 
  signal blk00000003_sig0000078d : STD_LOGIC; 
  signal blk00000003_sig0000078c : STD_LOGIC; 
  signal blk00000003_sig0000078b : STD_LOGIC; 
  signal blk00000003_sig0000078a : STD_LOGIC; 
  signal blk00000003_sig00000789 : STD_LOGIC; 
  signal blk00000003_sig00000788 : STD_LOGIC; 
  signal blk00000003_sig00000787 : STD_LOGIC; 
  signal blk00000003_sig00000786 : STD_LOGIC; 
  signal blk00000003_sig00000785 : STD_LOGIC; 
  signal blk00000003_sig00000784 : STD_LOGIC; 
  signal blk00000003_sig00000783 : STD_LOGIC; 
  signal blk00000003_sig00000782 : STD_LOGIC; 
  signal blk00000003_sig00000781 : STD_LOGIC; 
  signal blk00000003_sig00000780 : STD_LOGIC; 
  signal blk00000003_sig0000077f : STD_LOGIC; 
  signal blk00000003_sig0000077e : STD_LOGIC; 
  signal blk00000003_sig0000077d : STD_LOGIC; 
  signal blk00000003_sig0000077c : STD_LOGIC; 
  signal blk00000003_sig0000077b : STD_LOGIC; 
  signal blk00000003_sig0000077a : STD_LOGIC; 
  signal blk00000003_sig00000779 : STD_LOGIC; 
  signal blk00000003_sig00000778 : STD_LOGIC; 
  signal blk00000003_sig00000777 : STD_LOGIC; 
  signal blk00000003_sig00000776 : STD_LOGIC; 
  signal blk00000003_sig00000775 : STD_LOGIC; 
  signal blk00000003_sig00000774 : STD_LOGIC; 
  signal blk00000003_sig00000773 : STD_LOGIC; 
  signal blk00000003_sig00000772 : STD_LOGIC; 
  signal blk00000003_sig00000771 : STD_LOGIC; 
  signal blk00000003_sig00000770 : STD_LOGIC; 
  signal blk00000003_sig0000076f : STD_LOGIC; 
  signal blk00000003_sig0000076e : STD_LOGIC; 
  signal blk00000003_sig0000076d : STD_LOGIC; 
  signal blk00000003_sig0000076c : STD_LOGIC; 
  signal blk00000003_sig0000076b : STD_LOGIC; 
  signal blk00000003_sig0000076a : STD_LOGIC; 
  signal blk00000003_sig00000769 : STD_LOGIC; 
  signal blk00000003_sig00000768 : STD_LOGIC; 
  signal blk00000003_sig00000767 : STD_LOGIC; 
  signal blk00000003_sig00000766 : STD_LOGIC; 
  signal blk00000003_sig00000765 : STD_LOGIC; 
  signal blk00000003_sig00000764 : STD_LOGIC; 
  signal blk00000003_sig00000763 : STD_LOGIC; 
  signal blk00000003_sig00000762 : STD_LOGIC; 
  signal blk00000003_sig00000761 : STD_LOGIC; 
  signal blk00000003_sig00000760 : STD_LOGIC; 
  signal blk00000003_sig0000075f : STD_LOGIC; 
  signal blk00000003_sig0000075e : STD_LOGIC; 
  signal blk00000003_sig0000075d : STD_LOGIC; 
  signal blk00000003_sig0000075c : STD_LOGIC; 
  signal blk00000003_sig0000075b : STD_LOGIC; 
  signal blk00000003_sig0000075a : STD_LOGIC; 
  signal blk00000003_sig00000759 : STD_LOGIC; 
  signal blk00000003_sig00000758 : STD_LOGIC; 
  signal blk00000003_sig00000757 : STD_LOGIC; 
  signal blk00000003_sig00000756 : STD_LOGIC; 
  signal blk00000003_sig00000755 : STD_LOGIC; 
  signal blk00000003_sig00000754 : STD_LOGIC; 
  signal blk00000003_sig00000753 : STD_LOGIC; 
  signal blk00000003_sig00000752 : STD_LOGIC; 
  signal blk00000003_sig00000751 : STD_LOGIC; 
  signal blk00000003_sig00000750 : STD_LOGIC; 
  signal blk00000003_sig0000074f : STD_LOGIC; 
  signal blk00000003_sig0000074e : STD_LOGIC; 
  signal blk00000003_sig0000074d : STD_LOGIC; 
  signal blk00000003_sig0000074c : STD_LOGIC; 
  signal blk00000003_sig0000074b : STD_LOGIC; 
  signal blk00000003_sig0000074a : STD_LOGIC; 
  signal blk00000003_sig00000749 : STD_LOGIC; 
  signal blk00000003_sig00000748 : STD_LOGIC; 
  signal blk00000003_sig00000747 : STD_LOGIC; 
  signal blk00000003_sig00000746 : STD_LOGIC; 
  signal blk00000003_sig00000745 : STD_LOGIC; 
  signal blk00000003_sig00000744 : STD_LOGIC; 
  signal blk00000003_sig00000743 : STD_LOGIC; 
  signal blk00000003_sig00000742 : STD_LOGIC; 
  signal blk00000003_sig00000741 : STD_LOGIC; 
  signal blk00000003_sig00000740 : STD_LOGIC; 
  signal blk00000003_sig0000073f : STD_LOGIC; 
  signal blk00000003_sig0000073e : STD_LOGIC; 
  signal blk00000003_sig0000073d : STD_LOGIC; 
  signal blk00000003_sig0000073c : STD_LOGIC; 
  signal blk00000003_sig0000073b : STD_LOGIC; 
  signal blk00000003_sig0000073a : STD_LOGIC; 
  signal blk00000003_sig00000739 : STD_LOGIC; 
  signal blk00000003_sig00000738 : STD_LOGIC; 
  signal blk00000003_sig00000737 : STD_LOGIC; 
  signal blk00000003_sig00000736 : STD_LOGIC; 
  signal blk00000003_sig00000735 : STD_LOGIC; 
  signal blk00000003_sig00000734 : STD_LOGIC; 
  signal blk00000003_sig00000733 : STD_LOGIC; 
  signal blk00000003_sig00000732 : STD_LOGIC; 
  signal blk00000003_sig00000731 : STD_LOGIC; 
  signal blk00000003_sig00000730 : STD_LOGIC; 
  signal blk00000003_sig0000072f : STD_LOGIC; 
  signal blk00000003_sig0000072e : STD_LOGIC; 
  signal blk00000003_sig0000072d : STD_LOGIC; 
  signal blk00000003_sig0000072c : STD_LOGIC; 
  signal blk00000003_sig0000072b : STD_LOGIC; 
  signal blk00000003_sig0000072a : STD_LOGIC; 
  signal blk00000003_sig00000729 : STD_LOGIC; 
  signal blk00000003_sig00000728 : STD_LOGIC; 
  signal blk00000003_sig00000727 : STD_LOGIC; 
  signal blk00000003_sig00000726 : STD_LOGIC; 
  signal blk00000003_sig00000725 : STD_LOGIC; 
  signal blk00000003_sig00000724 : STD_LOGIC; 
  signal blk00000003_sig00000723 : STD_LOGIC; 
  signal blk00000003_sig00000722 : STD_LOGIC; 
  signal blk00000003_sig00000721 : STD_LOGIC; 
  signal blk00000003_sig00000720 : STD_LOGIC; 
  signal blk00000003_sig0000071f : STD_LOGIC; 
  signal blk00000003_sig0000071e : STD_LOGIC; 
  signal blk00000003_sig0000071d : STD_LOGIC; 
  signal blk00000003_sig0000071c : STD_LOGIC; 
  signal blk00000003_sig0000071b : STD_LOGIC; 
  signal blk00000003_sig0000071a : STD_LOGIC; 
  signal blk00000003_sig00000719 : STD_LOGIC; 
  signal blk00000003_sig00000718 : STD_LOGIC; 
  signal blk00000003_sig00000717 : STD_LOGIC; 
  signal blk00000003_sig00000716 : STD_LOGIC; 
  signal blk00000003_sig00000715 : STD_LOGIC; 
  signal blk00000003_sig00000714 : STD_LOGIC; 
  signal blk00000003_sig00000713 : STD_LOGIC; 
  signal blk00000003_sig00000712 : STD_LOGIC; 
  signal blk00000003_sig00000711 : STD_LOGIC; 
  signal blk00000003_sig00000710 : STD_LOGIC; 
  signal blk00000003_sig0000070f : STD_LOGIC; 
  signal blk00000003_sig0000070e : STD_LOGIC; 
  signal blk00000003_sig0000070d : STD_LOGIC; 
  signal blk00000003_sig0000070c : STD_LOGIC; 
  signal blk00000003_sig0000070b : STD_LOGIC; 
  signal blk00000003_sig0000070a : STD_LOGIC; 
  signal blk00000003_sig00000709 : STD_LOGIC; 
  signal blk00000003_sig00000708 : STD_LOGIC; 
  signal blk00000003_sig00000707 : STD_LOGIC; 
  signal blk00000003_sig00000706 : STD_LOGIC; 
  signal blk00000003_sig00000705 : STD_LOGIC; 
  signal blk00000003_sig00000704 : STD_LOGIC; 
  signal blk00000003_sig00000703 : STD_LOGIC; 
  signal blk00000003_sig00000702 : STD_LOGIC; 
  signal blk00000003_sig00000701 : STD_LOGIC; 
  signal blk00000003_sig00000700 : STD_LOGIC; 
  signal blk00000003_sig000006ff : STD_LOGIC; 
  signal blk00000003_sig000006fe : STD_LOGIC; 
  signal blk00000003_sig000006fd : STD_LOGIC; 
  signal blk00000003_sig000006fc : STD_LOGIC; 
  signal blk00000003_sig000006fb : STD_LOGIC; 
  signal blk00000003_sig000006fa : STD_LOGIC; 
  signal blk00000003_sig000006f9 : STD_LOGIC; 
  signal blk00000003_sig000006f8 : STD_LOGIC; 
  signal blk00000003_sig000006f7 : STD_LOGIC; 
  signal blk00000003_sig000006f6 : STD_LOGIC; 
  signal blk00000003_sig000006f5 : STD_LOGIC; 
  signal blk00000003_sig000006f4 : STD_LOGIC; 
  signal blk00000003_sig000006f3 : STD_LOGIC; 
  signal blk00000003_sig000006f2 : STD_LOGIC; 
  signal blk00000003_sig000006f1 : STD_LOGIC; 
  signal blk00000003_sig000006f0 : STD_LOGIC; 
  signal blk00000003_sig000006ef : STD_LOGIC; 
  signal blk00000003_sig000006ee : STD_LOGIC; 
  signal blk00000003_sig000006ed : STD_LOGIC; 
  signal blk00000003_sig000006ec : STD_LOGIC; 
  signal blk00000003_sig000006eb : STD_LOGIC; 
  signal blk00000003_sig000006ea : STD_LOGIC; 
  signal blk00000003_sig000006e9 : STD_LOGIC; 
  signal blk00000003_sig000006e8 : STD_LOGIC; 
  signal blk00000003_sig000006e7 : STD_LOGIC; 
  signal blk00000003_sig000006e6 : STD_LOGIC; 
  signal blk00000003_sig000006e5 : STD_LOGIC; 
  signal blk00000003_sig000006e4 : STD_LOGIC; 
  signal blk00000003_sig000006e3 : STD_LOGIC; 
  signal blk00000003_sig000006e2 : STD_LOGIC; 
  signal blk00000003_sig000006e1 : STD_LOGIC; 
  signal blk00000003_sig000006e0 : STD_LOGIC; 
  signal blk00000003_sig000006df : STD_LOGIC; 
  signal blk00000003_sig000006de : STD_LOGIC; 
  signal blk00000003_sig000006dd : STD_LOGIC; 
  signal blk00000003_sig000006dc : STD_LOGIC; 
  signal blk00000003_sig000006db : STD_LOGIC; 
  signal blk00000003_sig000006da : STD_LOGIC; 
  signal blk00000003_sig000006d9 : STD_LOGIC; 
  signal blk00000003_sig000006d8 : STD_LOGIC; 
  signal blk00000003_sig000006d7 : STD_LOGIC; 
  signal blk00000003_sig000006d6 : STD_LOGIC; 
  signal blk00000003_sig000006d5 : STD_LOGIC; 
  signal blk00000003_sig000006d4 : STD_LOGIC; 
  signal blk00000003_sig000006d3 : STD_LOGIC; 
  signal blk00000003_sig000006d2 : STD_LOGIC; 
  signal blk00000003_sig000006d1 : STD_LOGIC; 
  signal blk00000003_sig000006d0 : STD_LOGIC; 
  signal blk00000003_sig000006cf : STD_LOGIC; 
  signal blk00000003_sig000006ce : STD_LOGIC; 
  signal blk00000003_sig000006cd : STD_LOGIC; 
  signal blk00000003_sig000006cc : STD_LOGIC; 
  signal blk00000003_sig000006cb : STD_LOGIC; 
  signal blk00000003_sig000006ca : STD_LOGIC; 
  signal blk00000003_sig000006c9 : STD_LOGIC; 
  signal blk00000003_sig000006c8 : STD_LOGIC; 
  signal blk00000003_sig000006c7 : STD_LOGIC; 
  signal blk00000003_sig000006c6 : STD_LOGIC; 
  signal blk00000003_sig000006c5 : STD_LOGIC; 
  signal blk00000003_sig000006c4 : STD_LOGIC; 
  signal blk00000003_sig000006c3 : STD_LOGIC; 
  signal blk00000003_sig000006c2 : STD_LOGIC; 
  signal blk00000003_sig000006c1 : STD_LOGIC; 
  signal blk00000003_sig000006c0 : STD_LOGIC; 
  signal blk00000003_sig000006bf : STD_LOGIC; 
  signal blk00000003_sig000006be : STD_LOGIC; 
  signal blk00000003_sig000006bd : STD_LOGIC; 
  signal blk00000003_sig000006bc : STD_LOGIC; 
  signal blk00000003_sig000006bb : STD_LOGIC; 
  signal blk00000003_sig000006ba : STD_LOGIC; 
  signal blk00000003_sig000006b9 : STD_LOGIC; 
  signal blk00000003_sig000006b8 : STD_LOGIC; 
  signal blk00000003_sig000006b7 : STD_LOGIC; 
  signal blk00000003_sig000006b6 : STD_LOGIC; 
  signal blk00000003_sig000006b5 : STD_LOGIC; 
  signal blk00000003_sig000006b4 : STD_LOGIC; 
  signal blk00000003_sig000006b3 : STD_LOGIC; 
  signal blk00000003_sig000006b2 : STD_LOGIC; 
  signal blk00000003_sig000006b1 : STD_LOGIC; 
  signal blk00000003_sig000006b0 : STD_LOGIC; 
  signal blk00000003_sig000006af : STD_LOGIC; 
  signal blk00000003_sig000006ae : STD_LOGIC; 
  signal blk00000003_sig000006ad : STD_LOGIC; 
  signal blk00000003_sig000006ac : STD_LOGIC; 
  signal blk00000003_sig000006ab : STD_LOGIC; 
  signal blk00000003_sig000006aa : STD_LOGIC; 
  signal blk00000003_sig000006a9 : STD_LOGIC; 
  signal blk00000003_sig000006a8 : STD_LOGIC; 
  signal blk00000003_sig000006a7 : STD_LOGIC; 
  signal blk00000003_sig000006a6 : STD_LOGIC; 
  signal blk00000003_sig000006a5 : STD_LOGIC; 
  signal blk00000003_sig000006a4 : STD_LOGIC; 
  signal blk00000003_sig000006a3 : STD_LOGIC; 
  signal blk00000003_sig000006a2 : STD_LOGIC; 
  signal blk00000003_sig000006a1 : STD_LOGIC; 
  signal blk00000003_sig000006a0 : STD_LOGIC; 
  signal blk00000003_sig0000069f : STD_LOGIC; 
  signal blk00000003_sig0000069e : STD_LOGIC; 
  signal blk00000003_sig0000069d : STD_LOGIC; 
  signal blk00000003_sig0000069c : STD_LOGIC; 
  signal blk00000003_sig0000069b : STD_LOGIC; 
  signal blk00000003_sig0000069a : STD_LOGIC; 
  signal blk00000003_sig00000699 : STD_LOGIC; 
  signal blk00000003_sig00000698 : STD_LOGIC; 
  signal blk00000003_sig00000697 : STD_LOGIC; 
  signal blk00000003_sig00000696 : STD_LOGIC; 
  signal blk00000003_sig00000695 : STD_LOGIC; 
  signal blk00000003_sig00000694 : STD_LOGIC; 
  signal blk00000003_sig00000693 : STD_LOGIC; 
  signal blk00000003_sig00000692 : STD_LOGIC; 
  signal blk00000003_sig00000691 : STD_LOGIC; 
  signal blk00000003_sig00000690 : STD_LOGIC; 
  signal blk00000003_sig0000068f : STD_LOGIC; 
  signal blk00000003_sig0000068e : STD_LOGIC; 
  signal blk00000003_sig0000068d : STD_LOGIC; 
  signal blk00000003_sig0000068c : STD_LOGIC; 
  signal blk00000003_sig0000068b : STD_LOGIC; 
  signal blk00000003_sig0000068a : STD_LOGIC; 
  signal blk00000003_sig00000689 : STD_LOGIC; 
  signal blk00000003_sig00000688 : STD_LOGIC; 
  signal blk00000003_sig00000687 : STD_LOGIC; 
  signal blk00000003_sig00000686 : STD_LOGIC; 
  signal blk00000003_sig00000685 : STD_LOGIC; 
  signal blk00000003_sig00000684 : STD_LOGIC; 
  signal blk00000003_sig00000683 : STD_LOGIC; 
  signal blk00000003_sig00000682 : STD_LOGIC; 
  signal blk00000003_sig00000681 : STD_LOGIC; 
  signal blk00000003_sig00000680 : STD_LOGIC; 
  signal blk00000003_sig0000067f : STD_LOGIC; 
  signal blk00000003_sig0000067e : STD_LOGIC; 
  signal blk00000003_sig0000067d : STD_LOGIC; 
  signal blk00000003_sig0000067c : STD_LOGIC; 
  signal blk00000003_sig0000067b : STD_LOGIC; 
  signal blk00000003_sig0000067a : STD_LOGIC; 
  signal blk00000003_sig00000679 : STD_LOGIC; 
  signal blk00000003_sig00000678 : STD_LOGIC; 
  signal blk00000003_sig00000677 : STD_LOGIC; 
  signal blk00000003_sig00000676 : STD_LOGIC; 
  signal blk00000003_sig00000675 : STD_LOGIC; 
  signal blk00000003_sig00000674 : STD_LOGIC; 
  signal blk00000003_sig00000673 : STD_LOGIC; 
  signal blk00000003_sig00000672 : STD_LOGIC; 
  signal blk00000003_sig00000671 : STD_LOGIC; 
  signal blk00000003_sig00000670 : STD_LOGIC; 
  signal blk00000003_sig0000066f : STD_LOGIC; 
  signal blk00000003_sig0000066e : STD_LOGIC; 
  signal blk00000003_sig0000066d : STD_LOGIC; 
  signal blk00000003_sig0000066c : STD_LOGIC; 
  signal blk00000003_sig0000066b : STD_LOGIC; 
  signal blk00000003_sig0000066a : STD_LOGIC; 
  signal blk00000003_sig00000669 : STD_LOGIC; 
  signal blk00000003_sig00000668 : STD_LOGIC; 
  signal blk00000003_sig00000667 : STD_LOGIC; 
  signal blk00000003_sig00000666 : STD_LOGIC; 
  signal blk00000003_sig00000665 : STD_LOGIC; 
  signal blk00000003_sig00000664 : STD_LOGIC; 
  signal blk00000003_sig00000663 : STD_LOGIC; 
  signal blk00000003_sig00000662 : STD_LOGIC; 
  signal blk00000003_sig00000661 : STD_LOGIC; 
  signal blk00000003_sig00000660 : STD_LOGIC; 
  signal blk00000003_sig0000065f : STD_LOGIC; 
  signal blk00000003_sig0000065e : STD_LOGIC; 
  signal blk00000003_sig0000065d : STD_LOGIC; 
  signal blk00000003_sig0000065c : STD_LOGIC; 
  signal blk00000003_sig0000065b : STD_LOGIC; 
  signal blk00000003_sig0000065a : STD_LOGIC; 
  signal blk00000003_sig00000659 : STD_LOGIC; 
  signal blk00000003_sig00000658 : STD_LOGIC; 
  signal blk00000003_sig00000657 : STD_LOGIC; 
  signal blk00000003_sig00000656 : STD_LOGIC; 
  signal blk00000003_sig00000655 : STD_LOGIC; 
  signal blk00000003_sig00000654 : STD_LOGIC; 
  signal blk00000003_sig00000653 : STD_LOGIC; 
  signal blk00000003_sig00000652 : STD_LOGIC; 
  signal blk00000003_sig00000651 : STD_LOGIC; 
  signal blk00000003_sig00000650 : STD_LOGIC; 
  signal blk00000003_sig0000064f : STD_LOGIC; 
  signal blk00000003_sig0000064e : STD_LOGIC; 
  signal blk00000003_sig0000064d : STD_LOGIC; 
  signal blk00000003_sig0000064c : STD_LOGIC; 
  signal blk00000003_sig0000064b : STD_LOGIC; 
  signal blk00000003_sig0000064a : STD_LOGIC; 
  signal blk00000003_sig00000649 : STD_LOGIC; 
  signal blk00000003_sig00000648 : STD_LOGIC; 
  signal blk00000003_sig00000647 : STD_LOGIC; 
  signal blk00000003_sig00000646 : STD_LOGIC; 
  signal blk00000003_sig00000645 : STD_LOGIC; 
  signal blk00000003_sig00000644 : STD_LOGIC; 
  signal blk00000003_sig00000643 : STD_LOGIC; 
  signal blk00000003_sig00000642 : STD_LOGIC; 
  signal blk00000003_sig00000641 : STD_LOGIC; 
  signal blk00000003_sig00000640 : STD_LOGIC; 
  signal blk00000003_sig0000063f : STD_LOGIC; 
  signal blk00000003_sig0000063e : STD_LOGIC; 
  signal blk00000003_sig0000063d : STD_LOGIC; 
  signal blk00000003_sig0000063c : STD_LOGIC; 
  signal blk00000003_sig0000063b : STD_LOGIC; 
  signal blk00000003_sig0000063a : STD_LOGIC; 
  signal blk00000003_sig00000639 : STD_LOGIC; 
  signal blk00000003_sig00000638 : STD_LOGIC; 
  signal blk00000003_sig00000637 : STD_LOGIC; 
  signal blk00000003_sig00000636 : STD_LOGIC; 
  signal blk00000003_sig00000635 : STD_LOGIC; 
  signal blk00000003_sig00000634 : STD_LOGIC; 
  signal blk00000003_sig00000633 : STD_LOGIC; 
  signal blk00000003_sig00000632 : STD_LOGIC; 
  signal blk00000003_sig00000631 : STD_LOGIC; 
  signal blk00000003_sig00000630 : STD_LOGIC; 
  signal blk00000003_sig0000062f : STD_LOGIC; 
  signal blk00000003_sig0000062e : STD_LOGIC; 
  signal blk00000003_sig0000062d : STD_LOGIC; 
  signal blk00000003_sig0000062c : STD_LOGIC; 
  signal blk00000003_sig0000062b : STD_LOGIC; 
  signal blk00000003_sig0000062a : STD_LOGIC; 
  signal blk00000003_sig00000629 : STD_LOGIC; 
  signal blk00000003_sig00000628 : STD_LOGIC; 
  signal blk00000003_sig00000627 : STD_LOGIC; 
  signal blk00000003_sig00000626 : STD_LOGIC; 
  signal blk00000003_sig00000625 : STD_LOGIC; 
  signal blk00000003_sig00000624 : STD_LOGIC; 
  signal blk00000003_sig00000623 : STD_LOGIC; 
  signal blk00000003_sig00000622 : STD_LOGIC; 
  signal blk00000003_sig00000621 : STD_LOGIC; 
  signal blk00000003_sig00000620 : STD_LOGIC; 
  signal blk00000003_sig0000061f : STD_LOGIC; 
  signal blk00000003_sig0000061e : STD_LOGIC; 
  signal blk00000003_sig0000061d : STD_LOGIC; 
  signal blk00000003_sig0000061c : STD_LOGIC; 
  signal blk00000003_sig0000061b : STD_LOGIC; 
  signal blk00000003_sig0000061a : STD_LOGIC; 
  signal blk00000003_sig00000619 : STD_LOGIC; 
  signal blk00000003_sig00000618 : STD_LOGIC; 
  signal blk00000003_sig00000617 : STD_LOGIC; 
  signal blk00000003_sig00000616 : STD_LOGIC; 
  signal blk00000003_sig00000615 : STD_LOGIC; 
  signal blk00000003_sig00000614 : STD_LOGIC; 
  signal blk00000003_sig00000613 : STD_LOGIC; 
  signal blk00000003_sig00000612 : STD_LOGIC; 
  signal blk00000003_sig00000611 : STD_LOGIC; 
  signal blk00000003_sig00000610 : STD_LOGIC; 
  signal blk00000003_sig0000060f : STD_LOGIC; 
  signal blk00000003_sig0000060e : STD_LOGIC; 
  signal blk00000003_sig0000060d : STD_LOGIC; 
  signal blk00000003_sig0000060c : STD_LOGIC; 
  signal blk00000003_sig0000060b : STD_LOGIC; 
  signal blk00000003_sig0000060a : STD_LOGIC; 
  signal blk00000003_sig00000609 : STD_LOGIC; 
  signal blk00000003_sig00000608 : STD_LOGIC; 
  signal blk00000003_sig00000607 : STD_LOGIC; 
  signal blk00000003_sig00000606 : STD_LOGIC; 
  signal blk00000003_sig00000605 : STD_LOGIC; 
  signal blk00000003_sig00000604 : STD_LOGIC; 
  signal blk00000003_sig00000603 : STD_LOGIC; 
  signal blk00000003_sig00000602 : STD_LOGIC; 
  signal blk00000003_sig00000601 : STD_LOGIC; 
  signal blk00000003_sig00000600 : STD_LOGIC; 
  signal blk00000003_sig000005ff : STD_LOGIC; 
  signal blk00000003_sig000005fe : STD_LOGIC; 
  signal blk00000003_sig000005fd : STD_LOGIC; 
  signal blk00000003_sig000005fc : STD_LOGIC; 
  signal blk00000003_sig000005fb : STD_LOGIC; 
  signal blk00000003_sig000005fa : STD_LOGIC; 
  signal blk00000003_sig000005f9 : STD_LOGIC; 
  signal blk00000003_sig000005f8 : STD_LOGIC; 
  signal blk00000003_sig000005f7 : STD_LOGIC; 
  signal blk00000003_sig000005f6 : STD_LOGIC; 
  signal blk00000003_sig000005f5 : STD_LOGIC; 
  signal blk00000003_sig000005f4 : STD_LOGIC; 
  signal blk00000003_sig000005f3 : STD_LOGIC; 
  signal blk00000003_sig000005f2 : STD_LOGIC; 
  signal blk00000003_sig000005f1 : STD_LOGIC; 
  signal blk00000003_sig000005f0 : STD_LOGIC; 
  signal blk00000003_sig000005ef : STD_LOGIC; 
  signal blk00000003_sig000005ee : STD_LOGIC; 
  signal blk00000003_sig000005ed : STD_LOGIC; 
  signal blk00000003_sig000005ec : STD_LOGIC; 
  signal blk00000003_sig000005eb : STD_LOGIC; 
  signal blk00000003_sig000005ea : STD_LOGIC; 
  signal blk00000003_sig000005e9 : STD_LOGIC; 
  signal blk00000003_sig000005e8 : STD_LOGIC; 
  signal blk00000003_sig000005e7 : STD_LOGIC; 
  signal blk00000003_sig000005e6 : STD_LOGIC; 
  signal blk00000003_sig000005e5 : STD_LOGIC; 
  signal blk00000003_sig000005e4 : STD_LOGIC; 
  signal blk00000003_sig000005e3 : STD_LOGIC; 
  signal blk00000003_sig000005e2 : STD_LOGIC; 
  signal blk00000003_sig000005e1 : STD_LOGIC; 
  signal blk00000003_sig000005e0 : STD_LOGIC; 
  signal blk00000003_sig000005df : STD_LOGIC; 
  signal blk00000003_sig000005de : STD_LOGIC; 
  signal blk00000003_sig000005dd : STD_LOGIC; 
  signal blk00000003_sig000005dc : STD_LOGIC; 
  signal blk00000003_sig000005db : STD_LOGIC; 
  signal blk00000003_sig000005da : STD_LOGIC; 
  signal blk00000003_sig000005d9 : STD_LOGIC; 
  signal blk00000003_sig000005d8 : STD_LOGIC; 
  signal blk00000003_sig000005d7 : STD_LOGIC; 
  signal blk00000003_sig000005d6 : STD_LOGIC; 
  signal blk00000003_sig000005d5 : STD_LOGIC; 
  signal blk00000003_sig000005d4 : STD_LOGIC; 
  signal blk00000003_sig000005d3 : STD_LOGIC; 
  signal blk00000003_sig000005d2 : STD_LOGIC; 
  signal blk00000003_sig000005d1 : STD_LOGIC; 
  signal blk00000003_sig000005d0 : STD_LOGIC; 
  signal blk00000003_sig000005cf : STD_LOGIC; 
  signal blk00000003_sig000005ce : STD_LOGIC; 
  signal blk00000003_sig000005cd : STD_LOGIC; 
  signal blk00000003_sig000005cc : STD_LOGIC; 
  signal blk00000003_sig000005cb : STD_LOGIC; 
  signal blk00000003_sig000005ca : STD_LOGIC; 
  signal blk00000003_sig000005c9 : STD_LOGIC; 
  signal blk00000003_sig000005c8 : STD_LOGIC; 
  signal blk00000003_sig000005c7 : STD_LOGIC; 
  signal blk00000003_sig000005c6 : STD_LOGIC; 
  signal blk00000003_sig000005c5 : STD_LOGIC; 
  signal blk00000003_sig000005c4 : STD_LOGIC; 
  signal blk00000003_sig000005c3 : STD_LOGIC; 
  signal blk00000003_sig000005c2 : STD_LOGIC; 
  signal blk00000003_sig000005c1 : STD_LOGIC; 
  signal blk00000003_sig000005c0 : STD_LOGIC; 
  signal blk00000003_sig000005bf : STD_LOGIC; 
  signal blk00000003_sig000005be : STD_LOGIC; 
  signal blk00000003_sig000005bd : STD_LOGIC; 
  signal blk00000003_sig000005bc : STD_LOGIC; 
  signal blk00000003_sig000005bb : STD_LOGIC; 
  signal blk00000003_sig000005ba : STD_LOGIC; 
  signal blk00000003_sig000005b9 : STD_LOGIC; 
  signal blk00000003_sig000005b8 : STD_LOGIC; 
  signal blk00000003_sig000005b7 : STD_LOGIC; 
  signal blk00000003_sig000005b6 : STD_LOGIC; 
  signal blk00000003_sig000005b5 : STD_LOGIC; 
  signal blk00000003_sig000005b4 : STD_LOGIC; 
  signal blk00000003_sig000005b3 : STD_LOGIC; 
  signal blk00000003_sig000005b2 : STD_LOGIC; 
  signal blk00000003_sig000005b1 : STD_LOGIC; 
  signal blk00000003_sig000005b0 : STD_LOGIC; 
  signal blk00000003_sig000005af : STD_LOGIC; 
  signal blk00000003_sig000005ae : STD_LOGIC; 
  signal blk00000003_sig000005ad : STD_LOGIC; 
  signal blk00000003_sig000005ac : STD_LOGIC; 
  signal blk00000003_sig000005ab : STD_LOGIC; 
  signal blk00000003_sig000005aa : STD_LOGIC; 
  signal blk00000003_sig000005a9 : STD_LOGIC; 
  signal blk00000003_sig000005a8 : STD_LOGIC; 
  signal blk00000003_sig000005a7 : STD_LOGIC; 
  signal blk00000003_sig000005a6 : STD_LOGIC; 
  signal blk00000003_sig000005a5 : STD_LOGIC; 
  signal blk00000003_sig000005a4 : STD_LOGIC; 
  signal blk00000003_sig000005a3 : STD_LOGIC; 
  signal blk00000003_sig000005a2 : STD_LOGIC; 
  signal blk00000003_sig000005a1 : STD_LOGIC; 
  signal blk00000003_sig000005a0 : STD_LOGIC; 
  signal blk00000003_sig0000059f : STD_LOGIC; 
  signal blk00000003_sig0000059e : STD_LOGIC; 
  signal blk00000003_sig0000059d : STD_LOGIC; 
  signal blk00000003_sig0000059c : STD_LOGIC; 
  signal blk00000003_sig0000059b : STD_LOGIC; 
  signal blk00000003_sig0000059a : STD_LOGIC; 
  signal blk00000003_sig00000599 : STD_LOGIC; 
  signal blk00000003_sig00000598 : STD_LOGIC; 
  signal blk00000003_sig00000597 : STD_LOGIC; 
  signal blk00000003_sig00000596 : STD_LOGIC; 
  signal blk00000003_sig00000595 : STD_LOGIC; 
  signal blk00000003_sig00000594 : STD_LOGIC; 
  signal blk00000003_sig00000593 : STD_LOGIC; 
  signal blk00000003_sig00000592 : STD_LOGIC; 
  signal blk00000003_sig00000591 : STD_LOGIC; 
  signal blk00000003_sig00000590 : STD_LOGIC; 
  signal blk00000003_sig0000058f : STD_LOGIC; 
  signal blk00000003_sig0000058e : STD_LOGIC; 
  signal blk00000003_sig0000058d : STD_LOGIC; 
  signal blk00000003_sig0000058c : STD_LOGIC; 
  signal blk00000003_sig0000058b : STD_LOGIC; 
  signal blk00000003_sig0000058a : STD_LOGIC; 
  signal blk00000003_sig00000589 : STD_LOGIC; 
  signal blk00000003_sig00000588 : STD_LOGIC; 
  signal blk00000003_sig00000587 : STD_LOGIC; 
  signal blk00000003_sig00000586 : STD_LOGIC; 
  signal blk00000003_sig00000585 : STD_LOGIC; 
  signal blk00000003_sig00000584 : STD_LOGIC; 
  signal blk00000003_sig00000583 : STD_LOGIC; 
  signal blk00000003_sig00000582 : STD_LOGIC; 
  signal blk00000003_sig00000581 : STD_LOGIC; 
  signal blk00000003_sig00000580 : STD_LOGIC; 
  signal blk00000003_sig0000057f : STD_LOGIC; 
  signal blk00000003_sig0000057e : STD_LOGIC; 
  signal blk00000003_sig0000057d : STD_LOGIC; 
  signal blk00000003_sig0000057c : STD_LOGIC; 
  signal blk00000003_sig0000057b : STD_LOGIC; 
  signal blk00000003_sig0000057a : STD_LOGIC; 
  signal blk00000003_sig00000579 : STD_LOGIC; 
  signal blk00000003_sig00000578 : STD_LOGIC; 
  signal blk00000003_sig00000577 : STD_LOGIC; 
  signal blk00000003_sig00000576 : STD_LOGIC; 
  signal blk00000003_sig00000575 : STD_LOGIC; 
  signal blk00000003_sig00000574 : STD_LOGIC; 
  signal blk00000003_sig00000573 : STD_LOGIC; 
  signal blk00000003_sig00000572 : STD_LOGIC; 
  signal blk00000003_sig00000571 : STD_LOGIC; 
  signal blk00000003_sig00000570 : STD_LOGIC; 
  signal blk00000003_sig0000056f : STD_LOGIC; 
  signal blk00000003_sig0000056e : STD_LOGIC; 
  signal blk00000003_sig0000056d : STD_LOGIC; 
  signal blk00000003_sig0000056c : STD_LOGIC; 
  signal blk00000003_sig0000056b : STD_LOGIC; 
  signal blk00000003_sig0000056a : STD_LOGIC; 
  signal blk00000003_sig00000569 : STD_LOGIC; 
  signal blk00000003_sig00000568 : STD_LOGIC; 
  signal blk00000003_sig00000567 : STD_LOGIC; 
  signal blk00000003_sig00000566 : STD_LOGIC; 
  signal blk00000003_sig00000565 : STD_LOGIC; 
  signal blk00000003_sig00000564 : STD_LOGIC; 
  signal blk00000003_sig00000563 : STD_LOGIC; 
  signal blk00000003_sig00000562 : STD_LOGIC; 
  signal blk00000003_sig00000561 : STD_LOGIC; 
  signal blk00000003_sig00000560 : STD_LOGIC; 
  signal blk00000003_sig0000055f : STD_LOGIC; 
  signal blk00000003_sig0000055e : STD_LOGIC; 
  signal blk00000003_sig0000055d : STD_LOGIC; 
  signal blk00000003_sig0000055c : STD_LOGIC; 
  signal blk00000003_sig0000055b : STD_LOGIC; 
  signal blk00000003_sig0000055a : STD_LOGIC; 
  signal blk00000003_sig00000559 : STD_LOGIC; 
  signal blk00000003_sig00000558 : STD_LOGIC; 
  signal blk00000003_sig00000557 : STD_LOGIC; 
  signal blk00000003_sig00000556 : STD_LOGIC; 
  signal blk00000003_sig00000555 : STD_LOGIC; 
  signal blk00000003_sig00000554 : STD_LOGIC; 
  signal blk00000003_sig00000553 : STD_LOGIC; 
  signal blk00000003_sig00000552 : STD_LOGIC; 
  signal blk00000003_sig00000551 : STD_LOGIC; 
  signal blk00000003_sig00000550 : STD_LOGIC; 
  signal blk00000003_sig0000054f : STD_LOGIC; 
  signal blk00000003_sig0000054e : STD_LOGIC; 
  signal blk00000003_sig0000054d : STD_LOGIC; 
  signal blk00000003_sig0000054c : STD_LOGIC; 
  signal blk00000003_sig0000054b : STD_LOGIC; 
  signal blk00000003_sig0000054a : STD_LOGIC; 
  signal blk00000003_sig00000549 : STD_LOGIC; 
  signal blk00000003_sig00000548 : STD_LOGIC; 
  signal blk00000003_sig00000547 : STD_LOGIC; 
  signal blk00000003_sig00000546 : STD_LOGIC; 
  signal blk00000003_sig00000545 : STD_LOGIC; 
  signal blk00000003_sig00000544 : STD_LOGIC; 
  signal blk00000003_sig00000543 : STD_LOGIC; 
  signal blk00000003_sig00000542 : STD_LOGIC; 
  signal blk00000003_sig00000541 : STD_LOGIC; 
  signal blk00000003_sig00000540 : STD_LOGIC; 
  signal blk00000003_sig0000053f : STD_LOGIC; 
  signal blk00000003_sig0000053e : STD_LOGIC; 
  signal blk00000003_sig0000053d : STD_LOGIC; 
  signal blk00000003_sig0000053c : STD_LOGIC; 
  signal blk00000003_sig0000053b : STD_LOGIC; 
  signal blk00000003_sig0000053a : STD_LOGIC; 
  signal blk00000003_sig00000539 : STD_LOGIC; 
  signal blk00000003_sig00000538 : STD_LOGIC; 
  signal blk00000003_sig00000537 : STD_LOGIC; 
  signal blk00000003_sig00000536 : STD_LOGIC; 
  signal blk00000003_sig00000535 : STD_LOGIC; 
  signal blk00000003_sig00000534 : STD_LOGIC; 
  signal blk00000003_sig00000533 : STD_LOGIC; 
  signal blk00000003_sig00000532 : STD_LOGIC; 
  signal blk00000003_sig00000531 : STD_LOGIC; 
  signal blk00000003_sig00000530 : STD_LOGIC; 
  signal blk00000003_sig0000052f : STD_LOGIC; 
  signal blk00000003_sig0000052e : STD_LOGIC; 
  signal blk00000003_sig0000052d : STD_LOGIC; 
  signal blk00000003_sig0000052c : STD_LOGIC; 
  signal blk00000003_sig0000052b : STD_LOGIC; 
  signal blk00000003_sig0000052a : STD_LOGIC; 
  signal blk00000003_sig00000529 : STD_LOGIC; 
  signal blk00000003_sig00000528 : STD_LOGIC; 
  signal blk00000003_sig00000527 : STD_LOGIC; 
  signal blk00000003_sig00000526 : STD_LOGIC; 
  signal blk00000003_sig00000525 : STD_LOGIC; 
  signal blk00000003_sig00000524 : STD_LOGIC; 
  signal blk00000003_sig00000523 : STD_LOGIC; 
  signal blk00000003_sig00000522 : STD_LOGIC; 
  signal blk00000003_sig00000521 : STD_LOGIC; 
  signal blk00000003_sig00000520 : STD_LOGIC; 
  signal blk00000003_sig0000051f : STD_LOGIC; 
  signal blk00000003_sig0000051e : STD_LOGIC; 
  signal blk00000003_sig0000051d : STD_LOGIC; 
  signal blk00000003_sig0000051c : STD_LOGIC; 
  signal blk00000003_sig0000051b : STD_LOGIC; 
  signal blk00000003_sig0000051a : STD_LOGIC; 
  signal blk00000003_sig00000519 : STD_LOGIC; 
  signal blk00000003_sig00000518 : STD_LOGIC; 
  signal blk00000003_sig00000517 : STD_LOGIC; 
  signal blk00000003_sig00000516 : STD_LOGIC; 
  signal blk00000003_sig00000515 : STD_LOGIC; 
  signal blk00000003_sig00000514 : STD_LOGIC; 
  signal blk00000003_sig00000513 : STD_LOGIC; 
  signal blk00000003_sig00000512 : STD_LOGIC; 
  signal blk00000003_sig00000511 : STD_LOGIC; 
  signal blk00000003_sig00000510 : STD_LOGIC; 
  signal blk00000003_sig0000050f : STD_LOGIC; 
  signal blk00000003_sig0000050e : STD_LOGIC; 
  signal blk00000003_sig0000050d : STD_LOGIC; 
  signal blk00000003_sig0000050c : STD_LOGIC; 
  signal blk00000003_sig0000050b : STD_LOGIC; 
  signal blk00000003_sig0000050a : STD_LOGIC; 
  signal blk00000003_sig00000509 : STD_LOGIC; 
  signal blk00000003_sig00000508 : STD_LOGIC; 
  signal blk00000003_sig00000507 : STD_LOGIC; 
  signal blk00000003_sig00000506 : STD_LOGIC; 
  signal blk00000003_sig00000505 : STD_LOGIC; 
  signal blk00000003_sig00000504 : STD_LOGIC; 
  signal blk00000003_sig00000503 : STD_LOGIC; 
  signal blk00000003_sig00000502 : STD_LOGIC; 
  signal blk00000003_sig00000501 : STD_LOGIC; 
  signal blk00000003_sig00000500 : STD_LOGIC; 
  signal blk00000003_sig000004ff : STD_LOGIC; 
  signal blk00000003_sig000004fe : STD_LOGIC; 
  signal blk00000003_sig000004fd : STD_LOGIC; 
  signal blk00000003_sig000004fc : STD_LOGIC; 
  signal blk00000003_sig000004fb : STD_LOGIC; 
  signal blk00000003_sig000004fa : STD_LOGIC; 
  signal blk00000003_sig000004f9 : STD_LOGIC; 
  signal blk00000003_sig000004f8 : STD_LOGIC; 
  signal blk00000003_sig000004f7 : STD_LOGIC; 
  signal blk00000003_sig000004f6 : STD_LOGIC; 
  signal blk00000003_sig000004f5 : STD_LOGIC; 
  signal blk00000003_sig000004f4 : STD_LOGIC; 
  signal blk00000003_sig000004f3 : STD_LOGIC; 
  signal blk00000003_sig000004f2 : STD_LOGIC; 
  signal blk00000003_sig000004f1 : STD_LOGIC; 
  signal blk00000003_sig000004f0 : STD_LOGIC; 
  signal blk00000003_sig000004ef : STD_LOGIC; 
  signal blk00000003_sig000004ee : STD_LOGIC; 
  signal blk00000003_sig000004ed : STD_LOGIC; 
  signal blk00000003_sig000004ec : STD_LOGIC; 
  signal blk00000003_sig000004eb : STD_LOGIC; 
  signal blk00000003_sig000004ea : STD_LOGIC; 
  signal blk00000003_sig000004e9 : STD_LOGIC; 
  signal blk00000003_sig000004e8 : STD_LOGIC; 
  signal blk00000003_sig000004e7 : STD_LOGIC; 
  signal blk00000003_sig000004e6 : STD_LOGIC; 
  signal blk00000003_sig000004e5 : STD_LOGIC; 
  signal blk00000003_sig000004e4 : STD_LOGIC; 
  signal blk00000003_sig000004e3 : STD_LOGIC; 
  signal blk00000003_sig000004e2 : STD_LOGIC; 
  signal blk00000003_sig000004e1 : STD_LOGIC; 
  signal blk00000003_sig000004e0 : STD_LOGIC; 
  signal blk00000003_sig000004df : STD_LOGIC; 
  signal blk00000003_sig000004de : STD_LOGIC; 
  signal blk00000003_sig000004dd : STD_LOGIC; 
  signal blk00000003_sig000004dc : STD_LOGIC; 
  signal blk00000003_sig000004db : STD_LOGIC; 
  signal blk00000003_sig000004da : STD_LOGIC; 
  signal blk00000003_sig000004d9 : STD_LOGIC; 
  signal blk00000003_sig000004d8 : STD_LOGIC; 
  signal blk00000003_sig000004d7 : STD_LOGIC; 
  signal blk00000003_sig000004d6 : STD_LOGIC; 
  signal blk00000003_sig000004d5 : STD_LOGIC; 
  signal blk00000003_sig000004d4 : STD_LOGIC; 
  signal blk00000003_sig000004d3 : STD_LOGIC; 
  signal blk00000003_sig000004d2 : STD_LOGIC; 
  signal blk00000003_sig000004d1 : STD_LOGIC; 
  signal blk00000003_sig000004d0 : STD_LOGIC; 
  signal blk00000003_sig000004cf : STD_LOGIC; 
  signal blk00000003_sig000004ce : STD_LOGIC; 
  signal blk00000003_sig000004cd : STD_LOGIC; 
  signal blk00000003_sig000004cc : STD_LOGIC; 
  signal blk00000003_sig000004cb : STD_LOGIC; 
  signal blk00000003_sig000004ca : STD_LOGIC; 
  signal blk00000003_sig000004c9 : STD_LOGIC; 
  signal blk00000003_sig000004c8 : STD_LOGIC; 
  signal blk00000003_sig000004c7 : STD_LOGIC; 
  signal blk00000003_sig000004c6 : STD_LOGIC; 
  signal blk00000003_sig000004c5 : STD_LOGIC; 
  signal blk00000003_sig000004c4 : STD_LOGIC; 
  signal blk00000003_sig000004c3 : STD_LOGIC; 
  signal blk00000003_sig000004c2 : STD_LOGIC; 
  signal blk00000003_sig000004c1 : STD_LOGIC; 
  signal blk00000003_sig000004c0 : STD_LOGIC; 
  signal blk00000003_sig000004bf : STD_LOGIC; 
  signal blk00000003_sig000004be : STD_LOGIC; 
  signal blk00000003_sig000004bd : STD_LOGIC; 
  signal blk00000003_sig000004bc : STD_LOGIC; 
  signal blk00000003_sig000004bb : STD_LOGIC; 
  signal blk00000003_sig000004ba : STD_LOGIC; 
  signal blk00000003_sig000004b9 : STD_LOGIC; 
  signal blk00000003_sig000004b8 : STD_LOGIC; 
  signal blk00000003_sig000004b7 : STD_LOGIC; 
  signal blk00000003_sig000004b6 : STD_LOGIC; 
  signal blk00000003_sig000004b5 : STD_LOGIC; 
  signal blk00000003_sig000004b4 : STD_LOGIC; 
  signal blk00000003_sig000004b3 : STD_LOGIC; 
  signal blk00000003_sig000004b2 : STD_LOGIC; 
  signal blk00000003_sig000004b1 : STD_LOGIC; 
  signal blk00000003_sig000004b0 : STD_LOGIC; 
  signal blk00000003_sig000004af : STD_LOGIC; 
  signal blk00000003_sig000004ae : STD_LOGIC; 
  signal blk00000003_sig000004ad : STD_LOGIC; 
  signal blk00000003_sig000004ac : STD_LOGIC; 
  signal blk00000003_sig000004ab : STD_LOGIC; 
  signal blk00000003_sig000004aa : STD_LOGIC; 
  signal blk00000003_sig000004a9 : STD_LOGIC; 
  signal blk00000003_sig000004a8 : STD_LOGIC; 
  signal blk00000003_sig000004a7 : STD_LOGIC; 
  signal blk00000003_sig000004a6 : STD_LOGIC; 
  signal blk00000003_sig000004a5 : STD_LOGIC; 
  signal blk00000003_sig000004a4 : STD_LOGIC; 
  signal blk00000003_sig000004a3 : STD_LOGIC; 
  signal blk00000003_sig000004a2 : STD_LOGIC; 
  signal blk00000003_sig000004a1 : STD_LOGIC; 
  signal blk00000003_sig000004a0 : STD_LOGIC; 
  signal blk00000003_sig0000049f : STD_LOGIC; 
  signal blk00000003_sig0000049e : STD_LOGIC; 
  signal blk00000003_sig0000049d : STD_LOGIC; 
  signal blk00000003_sig0000049c : STD_LOGIC; 
  signal blk00000003_sig0000049b : STD_LOGIC; 
  signal blk00000003_sig0000049a : STD_LOGIC; 
  signal blk00000003_sig00000499 : STD_LOGIC; 
  signal blk00000003_sig00000498 : STD_LOGIC; 
  signal blk00000003_sig00000497 : STD_LOGIC; 
  signal blk00000003_sig00000496 : STD_LOGIC; 
  signal blk00000003_sig00000495 : STD_LOGIC; 
  signal blk00000003_sig00000494 : STD_LOGIC; 
  signal blk00000003_sig00000493 : STD_LOGIC; 
  signal blk00000003_sig00000492 : STD_LOGIC; 
  signal blk00000003_sig00000491 : STD_LOGIC; 
  signal blk00000003_sig00000490 : STD_LOGIC; 
  signal blk00000003_sig0000048f : STD_LOGIC; 
  signal blk00000003_sig0000048e : STD_LOGIC; 
  signal blk00000003_sig0000048d : STD_LOGIC; 
  signal blk00000003_sig0000048c : STD_LOGIC; 
  signal blk00000003_sig0000048b : STD_LOGIC; 
  signal blk00000003_sig0000048a : STD_LOGIC; 
  signal blk00000003_sig00000489 : STD_LOGIC; 
  signal blk00000003_sig00000488 : STD_LOGIC; 
  signal blk00000003_sig00000487 : STD_LOGIC; 
  signal blk00000003_sig00000486 : STD_LOGIC; 
  signal blk00000003_sig00000485 : STD_LOGIC; 
  signal blk00000003_sig00000484 : STD_LOGIC; 
  signal blk00000003_sig00000483 : STD_LOGIC; 
  signal blk00000003_sig00000482 : STD_LOGIC; 
  signal blk00000003_sig00000481 : STD_LOGIC; 
  signal blk00000003_sig00000480 : STD_LOGIC; 
  signal blk00000003_sig0000047f : STD_LOGIC; 
  signal blk00000003_sig0000047e : STD_LOGIC; 
  signal blk00000003_sig0000047d : STD_LOGIC; 
  signal blk00000003_sig0000047c : STD_LOGIC; 
  signal blk00000003_sig0000047b : STD_LOGIC; 
  signal blk00000003_sig0000047a : STD_LOGIC; 
  signal blk00000003_sig00000479 : STD_LOGIC; 
  signal blk00000003_sig00000478 : STD_LOGIC; 
  signal blk00000003_sig00000477 : STD_LOGIC; 
  signal blk00000003_sig00000476 : STD_LOGIC; 
  signal blk00000003_sig00000475 : STD_LOGIC; 
  signal blk00000003_sig00000474 : STD_LOGIC; 
  signal blk00000003_sig00000473 : STD_LOGIC; 
  signal blk00000003_sig00000472 : STD_LOGIC; 
  signal blk00000003_sig00000471 : STD_LOGIC; 
  signal blk00000003_sig00000470 : STD_LOGIC; 
  signal blk00000003_sig0000046f : STD_LOGIC; 
  signal blk00000003_sig0000046e : STD_LOGIC; 
  signal blk00000003_sig0000046d : STD_LOGIC; 
  signal blk00000003_sig0000046c : STD_LOGIC; 
  signal blk00000003_sig0000046b : STD_LOGIC; 
  signal blk00000003_sig0000046a : STD_LOGIC; 
  signal blk00000003_sig00000469 : STD_LOGIC; 
  signal blk00000003_sig00000468 : STD_LOGIC; 
  signal blk00000003_sig00000467 : STD_LOGIC; 
  signal blk00000003_sig00000466 : STD_LOGIC; 
  signal blk00000003_sig00000465 : STD_LOGIC; 
  signal blk00000003_sig00000464 : STD_LOGIC; 
  signal blk00000003_sig00000463 : STD_LOGIC; 
  signal blk00000003_sig00000462 : STD_LOGIC; 
  signal blk00000003_sig00000461 : STD_LOGIC; 
  signal blk00000003_sig00000460 : STD_LOGIC; 
  signal blk00000003_sig0000045f : STD_LOGIC; 
  signal blk00000003_sig0000045e : STD_LOGIC; 
  signal blk00000003_sig0000045d : STD_LOGIC; 
  signal blk00000003_sig0000045c : STD_LOGIC; 
  signal blk00000003_sig0000045b : STD_LOGIC; 
  signal blk00000003_sig0000045a : STD_LOGIC; 
  signal blk00000003_sig00000459 : STD_LOGIC; 
  signal blk00000003_sig00000458 : STD_LOGIC; 
  signal blk00000003_sig00000457 : STD_LOGIC; 
  signal blk00000003_sig00000456 : STD_LOGIC; 
  signal blk00000003_sig00000455 : STD_LOGIC; 
  signal blk00000003_sig00000454 : STD_LOGIC; 
  signal blk00000003_sig00000453 : STD_LOGIC; 
  signal blk00000003_sig00000452 : STD_LOGIC; 
  signal blk00000003_sig00000451 : STD_LOGIC; 
  signal blk00000003_sig00000450 : STD_LOGIC; 
  signal blk00000003_sig0000044f : STD_LOGIC; 
  signal blk00000003_sig0000044e : STD_LOGIC; 
  signal blk00000003_sig0000044d : STD_LOGIC; 
  signal blk00000003_sig0000044c : STD_LOGIC; 
  signal blk00000003_sig0000044b : STD_LOGIC; 
  signal blk00000003_sig0000044a : STD_LOGIC; 
  signal blk00000003_sig00000449 : STD_LOGIC; 
  signal blk00000003_sig00000448 : STD_LOGIC; 
  signal blk00000003_sig00000447 : STD_LOGIC; 
  signal blk00000003_sig00000446 : STD_LOGIC; 
  signal blk00000003_sig00000445 : STD_LOGIC; 
  signal blk00000003_sig00000444 : STD_LOGIC; 
  signal blk00000003_sig00000443 : STD_LOGIC; 
  signal blk00000003_sig00000442 : STD_LOGIC; 
  signal blk00000003_sig00000441 : STD_LOGIC; 
  signal blk00000003_sig00000440 : STD_LOGIC; 
  signal blk00000003_sig0000043f : STD_LOGIC; 
  signal blk00000003_sig0000043e : STD_LOGIC; 
  signal blk00000003_sig0000043d : STD_LOGIC; 
  signal blk00000003_sig0000043c : STD_LOGIC; 
  signal blk00000003_sig0000043b : STD_LOGIC; 
  signal blk00000003_sig0000043a : STD_LOGIC; 
  signal blk00000003_sig00000439 : STD_LOGIC; 
  signal blk00000003_sig00000438 : STD_LOGIC; 
  signal blk00000003_sig00000437 : STD_LOGIC; 
  signal blk00000003_sig00000436 : STD_LOGIC; 
  signal blk00000003_sig00000435 : STD_LOGIC; 
  signal blk00000003_sig00000434 : STD_LOGIC; 
  signal blk00000003_sig00000433 : STD_LOGIC; 
  signal blk00000003_sig00000432 : STD_LOGIC; 
  signal blk00000003_sig00000431 : STD_LOGIC; 
  signal blk00000003_sig00000430 : STD_LOGIC; 
  signal blk00000003_sig0000042f : STD_LOGIC; 
  signal blk00000003_sig0000042e : STD_LOGIC; 
  signal blk00000003_sig0000042d : STD_LOGIC; 
  signal blk00000003_sig0000042c : STD_LOGIC; 
  signal blk00000003_sig0000042b : STD_LOGIC; 
  signal blk00000003_sig0000042a : STD_LOGIC; 
  signal blk00000003_sig00000429 : STD_LOGIC; 
  signal blk00000003_sig00000428 : STD_LOGIC; 
  signal blk00000003_sig00000427 : STD_LOGIC; 
  signal blk00000003_sig00000426 : STD_LOGIC; 
  signal blk00000003_sig00000425 : STD_LOGIC; 
  signal blk00000003_sig00000424 : STD_LOGIC; 
  signal blk00000003_sig00000423 : STD_LOGIC; 
  signal blk00000003_sig00000422 : STD_LOGIC; 
  signal blk00000003_sig00000421 : STD_LOGIC; 
  signal blk00000003_sig00000420 : STD_LOGIC; 
  signal blk00000003_sig0000041f : STD_LOGIC; 
  signal blk00000003_sig0000041e : STD_LOGIC; 
  signal blk00000003_sig0000041d : STD_LOGIC; 
  signal blk00000003_sig0000041c : STD_LOGIC; 
  signal blk00000003_sig0000041b : STD_LOGIC; 
  signal blk00000003_sig0000041a : STD_LOGIC; 
  signal blk00000003_sig00000419 : STD_LOGIC; 
  signal blk00000003_sig00000418 : STD_LOGIC; 
  signal blk00000003_sig00000417 : STD_LOGIC; 
  signal blk00000003_sig00000416 : STD_LOGIC; 
  signal blk00000003_sig00000415 : STD_LOGIC; 
  signal blk00000003_sig00000414 : STD_LOGIC; 
  signal blk00000003_sig00000413 : STD_LOGIC; 
  signal blk00000003_sig00000412 : STD_LOGIC; 
  signal blk00000003_sig00000411 : STD_LOGIC; 
  signal blk00000003_sig00000410 : STD_LOGIC; 
  signal blk00000003_sig0000040f : STD_LOGIC; 
  signal blk00000003_sig0000040e : STD_LOGIC; 
  signal blk00000003_sig0000040d : STD_LOGIC; 
  signal blk00000003_sig0000040c : STD_LOGIC; 
  signal blk00000003_sig0000040b : STD_LOGIC; 
  signal blk00000003_sig0000040a : STD_LOGIC; 
  signal blk00000003_sig00000409 : STD_LOGIC; 
  signal blk00000003_sig00000408 : STD_LOGIC; 
  signal blk00000003_sig00000407 : STD_LOGIC; 
  signal blk00000003_sig00000406 : STD_LOGIC; 
  signal blk00000003_sig00000405 : STD_LOGIC; 
  signal blk00000003_sig00000404 : STD_LOGIC; 
  signal blk00000003_sig00000403 : STD_LOGIC; 
  signal blk00000003_sig00000402 : STD_LOGIC; 
  signal blk00000003_sig00000401 : STD_LOGIC; 
  signal blk00000003_sig00000400 : STD_LOGIC; 
  signal blk00000003_sig000003ff : STD_LOGIC; 
  signal blk00000003_sig000003fe : STD_LOGIC; 
  signal blk00000003_sig000003fd : STD_LOGIC; 
  signal blk00000003_sig000003fc : STD_LOGIC; 
  signal blk00000003_sig000003fb : STD_LOGIC; 
  signal blk00000003_sig000003fa : STD_LOGIC; 
  signal blk00000003_sig000003f9 : STD_LOGIC; 
  signal blk00000003_sig000003f8 : STD_LOGIC; 
  signal blk00000003_sig000003f7 : STD_LOGIC; 
  signal blk00000003_sig000003f6 : STD_LOGIC; 
  signal blk00000003_sig000003f5 : STD_LOGIC; 
  signal blk00000003_sig000003f4 : STD_LOGIC; 
  signal blk00000003_sig000003f3 : STD_LOGIC; 
  signal blk00000003_sig000003f2 : STD_LOGIC; 
  signal blk00000003_sig000003f1 : STD_LOGIC; 
  signal blk00000003_sig000003f0 : STD_LOGIC; 
  signal blk00000003_sig000003ef : STD_LOGIC; 
  signal blk00000003_sig000003ee : STD_LOGIC; 
  signal blk00000003_sig000003ed : STD_LOGIC; 
  signal blk00000003_sig000003ec : STD_LOGIC; 
  signal blk00000003_sig000003eb : STD_LOGIC; 
  signal blk00000003_sig000003ea : STD_LOGIC; 
  signal blk00000003_sig000003e9 : STD_LOGIC; 
  signal blk00000003_sig000003e8 : STD_LOGIC; 
  signal blk00000003_sig000003e7 : STD_LOGIC; 
  signal blk00000003_sig000003e6 : STD_LOGIC; 
  signal blk00000003_sig000003e5 : STD_LOGIC; 
  signal blk00000003_sig000003e4 : STD_LOGIC; 
  signal blk00000003_sig000003e3 : STD_LOGIC; 
  signal blk00000003_sig000003e2 : STD_LOGIC; 
  signal blk00000003_sig000003e1 : STD_LOGIC; 
  signal blk00000003_sig000003e0 : STD_LOGIC; 
  signal blk00000003_sig000003df : STD_LOGIC; 
  signal blk00000003_sig000003de : STD_LOGIC; 
  signal blk00000003_sig000003dd : STD_LOGIC; 
  signal blk00000003_sig000003dc : STD_LOGIC; 
  signal blk00000003_sig000003db : STD_LOGIC; 
  signal blk00000003_sig000003da : STD_LOGIC; 
  signal blk00000003_sig000003d9 : STD_LOGIC; 
  signal blk00000003_sig000003d8 : STD_LOGIC; 
  signal blk00000003_sig000003d7 : STD_LOGIC; 
  signal blk00000003_sig000003d6 : STD_LOGIC; 
  signal blk00000003_sig000003d5 : STD_LOGIC; 
  signal blk00000003_sig000003d4 : STD_LOGIC; 
  signal blk00000003_sig000003d3 : STD_LOGIC; 
  signal blk00000003_sig000003d2 : STD_LOGIC; 
  signal blk00000003_sig000003d1 : STD_LOGIC; 
  signal blk00000003_sig000003d0 : STD_LOGIC; 
  signal blk00000003_sig000003cf : STD_LOGIC; 
  signal blk00000003_sig000003ce : STD_LOGIC; 
  signal blk00000003_sig000003cd : STD_LOGIC; 
  signal blk00000003_sig000003cc : STD_LOGIC; 
  signal blk00000003_sig000003cb : STD_LOGIC; 
  signal blk00000003_sig000003ca : STD_LOGIC; 
  signal blk00000003_sig000003c9 : STD_LOGIC; 
  signal blk00000003_sig000003c8 : STD_LOGIC; 
  signal blk00000003_sig000003c7 : STD_LOGIC; 
  signal blk00000003_sig000003c6 : STD_LOGIC; 
  signal blk00000003_sig000003c5 : STD_LOGIC; 
  signal blk00000003_sig000003c4 : STD_LOGIC; 
  signal blk00000003_sig000003c3 : STD_LOGIC; 
  signal blk00000003_sig000003c2 : STD_LOGIC; 
  signal blk00000003_sig000003c1 : STD_LOGIC; 
  signal blk00000003_sig000003c0 : STD_LOGIC; 
  signal blk00000003_sig000003bf : STD_LOGIC; 
  signal blk00000003_sig000003be : STD_LOGIC; 
  signal blk00000003_sig000003bd : STD_LOGIC; 
  signal blk00000003_sig000003bc : STD_LOGIC; 
  signal blk00000003_sig000003bb : STD_LOGIC; 
  signal blk00000003_sig000003ba : STD_LOGIC; 
  signal blk00000003_sig000003b9 : STD_LOGIC; 
  signal blk00000003_sig000003b8 : STD_LOGIC; 
  signal blk00000003_sig000003b7 : STD_LOGIC; 
  signal blk00000003_sig000003b6 : STD_LOGIC; 
  signal blk00000003_sig000003b5 : STD_LOGIC; 
  signal blk00000003_sig000003b4 : STD_LOGIC; 
  signal blk00000003_sig000003b3 : STD_LOGIC; 
  signal blk00000003_sig000003b2 : STD_LOGIC; 
  signal blk00000003_sig000003b1 : STD_LOGIC; 
  signal blk00000003_sig000003b0 : STD_LOGIC; 
  signal blk00000003_sig000003af : STD_LOGIC; 
  signal blk00000003_sig000003ae : STD_LOGIC; 
  signal blk00000003_sig000003ad : STD_LOGIC; 
  signal blk00000003_sig000003ac : STD_LOGIC; 
  signal blk00000003_sig000003ab : STD_LOGIC; 
  signal blk00000003_sig000003aa : STD_LOGIC; 
  signal blk00000003_sig000003a9 : STD_LOGIC; 
  signal blk00000003_sig000003a8 : STD_LOGIC; 
  signal blk00000003_sig000003a7 : STD_LOGIC; 
  signal blk00000003_sig000003a6 : STD_LOGIC; 
  signal blk00000003_sig000003a5 : STD_LOGIC; 
  signal blk00000003_sig000003a4 : STD_LOGIC; 
  signal blk00000003_sig000003a3 : STD_LOGIC; 
  signal blk00000003_sig000003a2 : STD_LOGIC; 
  signal blk00000003_sig000003a1 : STD_LOGIC; 
  signal blk00000003_sig000003a0 : STD_LOGIC; 
  signal blk00000003_sig0000039f : STD_LOGIC; 
  signal blk00000003_sig0000039e : STD_LOGIC; 
  signal blk00000003_sig0000039d : STD_LOGIC; 
  signal blk00000003_sig0000039c : STD_LOGIC; 
  signal blk00000003_sig0000039b : STD_LOGIC; 
  signal blk00000003_sig0000039a : STD_LOGIC; 
  signal blk00000003_sig00000399 : STD_LOGIC; 
  signal blk00000003_sig00000398 : STD_LOGIC; 
  signal blk00000003_sig00000397 : STD_LOGIC; 
  signal blk00000003_sig00000396 : STD_LOGIC; 
  signal blk00000003_sig00000395 : STD_LOGIC; 
  signal blk00000003_sig00000394 : STD_LOGIC; 
  signal blk00000003_sig00000393 : STD_LOGIC; 
  signal blk00000003_sig00000392 : STD_LOGIC; 
  signal blk00000003_sig00000391 : STD_LOGIC; 
  signal blk00000003_sig00000390 : STD_LOGIC; 
  signal blk00000003_sig0000038f : STD_LOGIC; 
  signal blk00000003_sig0000038e : STD_LOGIC; 
  signal blk00000003_sig0000038d : STD_LOGIC; 
  signal blk00000003_sig0000038c : STD_LOGIC; 
  signal blk00000003_sig0000038b : STD_LOGIC; 
  signal blk00000003_sig0000038a : STD_LOGIC; 
  signal blk00000003_sig00000389 : STD_LOGIC; 
  signal blk00000003_sig00000388 : STD_LOGIC; 
  signal blk00000003_sig00000387 : STD_LOGIC; 
  signal blk00000003_sig00000386 : STD_LOGIC; 
  signal blk00000003_sig00000385 : STD_LOGIC; 
  signal blk00000003_sig00000384 : STD_LOGIC; 
  signal blk00000003_sig00000383 : STD_LOGIC; 
  signal blk00000003_sig00000382 : STD_LOGIC; 
  signal blk00000003_sig00000381 : STD_LOGIC; 
  signal blk00000003_sig00000380 : STD_LOGIC; 
  signal blk00000003_sig0000037f : STD_LOGIC; 
  signal blk00000003_sig0000037e : STD_LOGIC; 
  signal blk00000003_sig0000037d : STD_LOGIC; 
  signal blk00000003_sig0000037c : STD_LOGIC; 
  signal blk00000003_sig0000037b : STD_LOGIC; 
  signal blk00000003_sig0000037a : STD_LOGIC; 
  signal blk00000003_sig00000379 : STD_LOGIC; 
  signal blk00000003_sig00000378 : STD_LOGIC; 
  signal blk00000003_sig00000377 : STD_LOGIC; 
  signal blk00000003_sig00000376 : STD_LOGIC; 
  signal blk00000003_sig00000375 : STD_LOGIC; 
  signal blk00000003_sig00000374 : STD_LOGIC; 
  signal blk00000003_sig00000373 : STD_LOGIC; 
  signal blk00000003_sig00000372 : STD_LOGIC; 
  signal blk00000003_sig00000371 : STD_LOGIC; 
  signal blk00000003_sig00000370 : STD_LOGIC; 
  signal blk00000003_sig0000036f : STD_LOGIC; 
  signal blk00000003_sig0000036e : STD_LOGIC; 
  signal blk00000003_sig0000036d : STD_LOGIC; 
  signal blk00000003_sig0000036c : STD_LOGIC; 
  signal blk00000003_sig0000036b : STD_LOGIC; 
  signal blk00000003_sig0000036a : STD_LOGIC; 
  signal blk00000003_sig00000369 : STD_LOGIC; 
  signal blk00000003_sig00000368 : STD_LOGIC; 
  signal blk00000003_sig00000367 : STD_LOGIC; 
  signal blk00000003_sig00000366 : STD_LOGIC; 
  signal blk00000003_sig00000365 : STD_LOGIC; 
  signal blk00000003_sig00000364 : STD_LOGIC; 
  signal blk00000003_sig00000363 : STD_LOGIC; 
  signal blk00000003_sig00000362 : STD_LOGIC; 
  signal blk00000003_sig00000361 : STD_LOGIC; 
  signal blk00000003_sig00000360 : STD_LOGIC; 
  signal blk00000003_sig0000035f : STD_LOGIC; 
  signal blk00000003_sig0000035e : STD_LOGIC; 
  signal blk00000003_sig0000035d : STD_LOGIC; 
  signal blk00000003_sig0000035c : STD_LOGIC; 
  signal blk00000003_sig0000035b : STD_LOGIC; 
  signal blk00000003_sig0000035a : STD_LOGIC; 
  signal blk00000003_sig00000359 : STD_LOGIC; 
  signal blk00000003_sig00000358 : STD_LOGIC; 
  signal blk00000003_sig00000357 : STD_LOGIC; 
  signal blk00000003_sig00000356 : STD_LOGIC; 
  signal blk00000003_sig00000355 : STD_LOGIC; 
  signal blk00000003_sig00000354 : STD_LOGIC; 
  signal blk00000003_sig00000353 : STD_LOGIC; 
  signal blk00000003_sig00000352 : STD_LOGIC; 
  signal blk00000003_sig00000351 : STD_LOGIC; 
  signal blk00000003_sig00000350 : STD_LOGIC; 
  signal blk00000003_sig0000034f : STD_LOGIC; 
  signal blk00000003_sig0000034e : STD_LOGIC; 
  signal blk00000003_sig0000034d : STD_LOGIC; 
  signal blk00000003_sig0000034c : STD_LOGIC; 
  signal blk00000003_sig0000034b : STD_LOGIC; 
  signal blk00000003_sig0000034a : STD_LOGIC; 
  signal blk00000003_sig00000349 : STD_LOGIC; 
  signal blk00000003_sig00000348 : STD_LOGIC; 
  signal blk00000003_sig00000347 : STD_LOGIC; 
  signal blk00000003_sig00000346 : STD_LOGIC; 
  signal blk00000003_sig00000345 : STD_LOGIC; 
  signal blk00000003_sig00000344 : STD_LOGIC; 
  signal blk00000003_sig00000343 : STD_LOGIC; 
  signal blk00000003_sig00000342 : STD_LOGIC; 
  signal blk00000003_sig00000341 : STD_LOGIC; 
  signal blk00000003_sig00000340 : STD_LOGIC; 
  signal blk00000003_sig0000033f : STD_LOGIC; 
  signal blk00000003_sig0000033e : STD_LOGIC; 
  signal blk00000003_sig0000033d : STD_LOGIC; 
  signal blk00000003_sig0000033c : STD_LOGIC; 
  signal blk00000003_sig0000033b : STD_LOGIC; 
  signal blk00000003_sig0000033a : STD_LOGIC; 
  signal blk00000003_sig00000339 : STD_LOGIC; 
  signal blk00000003_sig00000338 : STD_LOGIC; 
  signal blk00000003_sig00000337 : STD_LOGIC; 
  signal blk00000003_sig00000336 : STD_LOGIC; 
  signal blk00000003_sig00000335 : STD_LOGIC; 
  signal blk00000003_sig00000334 : STD_LOGIC; 
  signal blk00000003_sig00000333 : STD_LOGIC; 
  signal blk00000003_sig00000332 : STD_LOGIC; 
  signal blk00000003_sig00000331 : STD_LOGIC; 
  signal blk00000003_sig00000330 : STD_LOGIC; 
  signal blk00000003_sig0000032f : STD_LOGIC; 
  signal blk00000003_sig0000032e : STD_LOGIC; 
  signal blk00000003_sig0000032d : STD_LOGIC; 
  signal blk00000003_sig0000032c : STD_LOGIC; 
  signal blk00000003_sig0000032b : STD_LOGIC; 
  signal blk00000003_sig0000032a : STD_LOGIC; 
  signal blk00000003_sig00000329 : STD_LOGIC; 
  signal blk00000003_sig00000328 : STD_LOGIC; 
  signal blk00000003_sig00000327 : STD_LOGIC; 
  signal blk00000003_sig00000326 : STD_LOGIC; 
  signal blk00000003_sig00000325 : STD_LOGIC; 
  signal blk00000003_sig00000324 : STD_LOGIC; 
  signal blk00000003_sig00000323 : STD_LOGIC; 
  signal blk00000003_sig00000322 : STD_LOGIC; 
  signal blk00000003_sig00000321 : STD_LOGIC; 
  signal blk00000003_sig00000320 : STD_LOGIC; 
  signal blk00000003_sig0000031f : STD_LOGIC; 
  signal blk00000003_sig0000031e : STD_LOGIC; 
  signal blk00000003_sig0000031d : STD_LOGIC; 
  signal blk00000003_sig0000031c : STD_LOGIC; 
  signal blk00000003_sig0000031b : STD_LOGIC; 
  signal blk00000003_sig0000031a : STD_LOGIC; 
  signal blk00000003_sig00000319 : STD_LOGIC; 
  signal blk00000003_sig00000318 : STD_LOGIC; 
  signal blk00000003_sig00000317 : STD_LOGIC; 
  signal blk00000003_sig00000316 : STD_LOGIC; 
  signal blk00000003_sig00000315 : STD_LOGIC; 
  signal blk00000003_sig00000314 : STD_LOGIC; 
  signal blk00000003_sig00000313 : STD_LOGIC; 
  signal blk00000003_sig00000312 : STD_LOGIC; 
  signal blk00000003_sig00000311 : STD_LOGIC; 
  signal blk00000003_sig00000310 : STD_LOGIC; 
  signal blk00000003_sig0000030f : STD_LOGIC; 
  signal blk00000003_sig0000030e : STD_LOGIC; 
  signal blk00000003_sig0000030d : STD_LOGIC; 
  signal blk00000003_sig0000030c : STD_LOGIC; 
  signal blk00000003_sig0000030b : STD_LOGIC; 
  signal blk00000003_sig0000030a : STD_LOGIC; 
  signal blk00000003_sig00000309 : STD_LOGIC; 
  signal blk00000003_sig00000308 : STD_LOGIC; 
  signal blk00000003_sig00000307 : STD_LOGIC; 
  signal blk00000003_sig00000306 : STD_LOGIC; 
  signal blk00000003_sig00000305 : STD_LOGIC; 
  signal blk00000003_sig00000304 : STD_LOGIC; 
  signal blk00000003_sig00000303 : STD_LOGIC; 
  signal blk00000003_sig00000302 : STD_LOGIC; 
  signal blk00000003_sig00000301 : STD_LOGIC; 
  signal blk00000003_sig00000300 : STD_LOGIC; 
  signal blk00000003_sig000002ff : STD_LOGIC; 
  signal blk00000003_sig000002fe : STD_LOGIC; 
  signal blk00000003_sig000002fd : STD_LOGIC; 
  signal blk00000003_sig000002fc : STD_LOGIC; 
  signal blk00000003_sig000002fb : STD_LOGIC; 
  signal blk00000003_sig000002fa : STD_LOGIC; 
  signal blk00000003_sig000002f9 : STD_LOGIC; 
  signal blk00000003_sig000002f8 : STD_LOGIC; 
  signal blk00000003_sig000002f7 : STD_LOGIC; 
  signal blk00000003_sig000002f6 : STD_LOGIC; 
  signal blk00000003_sig000002f5 : STD_LOGIC; 
  signal blk00000003_sig000002f4 : STD_LOGIC; 
  signal blk00000003_sig000002f3 : STD_LOGIC; 
  signal blk00000003_sig000002f2 : STD_LOGIC; 
  signal blk00000003_sig000002f1 : STD_LOGIC; 
  signal blk00000003_sig000002f0 : STD_LOGIC; 
  signal blk00000003_sig000002ef : STD_LOGIC; 
  signal blk00000003_sig000002ee : STD_LOGIC; 
  signal blk00000003_sig000002ed : STD_LOGIC; 
  signal blk00000003_sig000002ec : STD_LOGIC; 
  signal blk00000003_sig000002eb : STD_LOGIC; 
  signal blk00000003_sig000002ea : STD_LOGIC; 
  signal blk00000003_sig000002e9 : STD_LOGIC; 
  signal blk00000003_sig000002e8 : STD_LOGIC; 
  signal blk00000003_sig000002e7 : STD_LOGIC; 
  signal blk00000003_sig000002e6 : STD_LOGIC; 
  signal blk00000003_sig000002e5 : STD_LOGIC; 
  signal blk00000003_sig000002e4 : STD_LOGIC; 
  signal blk00000003_sig000002e3 : STD_LOGIC; 
  signal blk00000003_sig000002e2 : STD_LOGIC; 
  signal blk00000003_sig000002e1 : STD_LOGIC; 
  signal blk00000003_sig000002e0 : STD_LOGIC; 
  signal blk00000003_sig000002df : STD_LOGIC; 
  signal blk00000003_sig000002de : STD_LOGIC; 
  signal blk00000003_sig000002dd : STD_LOGIC; 
  signal blk00000003_sig000002dc : STD_LOGIC; 
  signal blk00000003_sig000002db : STD_LOGIC; 
  signal blk00000003_sig000002da : STD_LOGIC; 
  signal blk00000003_sig000002d9 : STD_LOGIC; 
  signal blk00000003_sig000002d8 : STD_LOGIC; 
  signal blk00000003_sig000002d7 : STD_LOGIC; 
  signal blk00000003_sig000002d6 : STD_LOGIC; 
  signal blk00000003_sig000002d5 : STD_LOGIC; 
  signal blk00000003_sig000002d4 : STD_LOGIC; 
  signal blk00000003_sig000002d3 : STD_LOGIC; 
  signal blk00000003_sig000002d2 : STD_LOGIC; 
  signal blk00000003_sig000002d1 : STD_LOGIC; 
  signal blk00000003_sig000002d0 : STD_LOGIC; 
  signal blk00000003_sig000002cf : STD_LOGIC; 
  signal blk00000003_sig000002ce : STD_LOGIC; 
  signal blk00000003_sig000002cd : STD_LOGIC; 
  signal blk00000003_sig000002cc : STD_LOGIC; 
  signal blk00000003_sig000002cb : STD_LOGIC; 
  signal blk00000003_sig000002ca : STD_LOGIC; 
  signal blk00000003_sig000002c9 : STD_LOGIC; 
  signal blk00000003_sig000002c8 : STD_LOGIC; 
  signal blk00000003_sig000002c7 : STD_LOGIC; 
  signal blk00000003_sig000002c6 : STD_LOGIC; 
  signal blk00000003_sig000002c5 : STD_LOGIC; 
  signal blk00000003_sig000002c4 : STD_LOGIC; 
  signal blk00000003_sig000002c3 : STD_LOGIC; 
  signal blk00000003_sig000002c2 : STD_LOGIC; 
  signal blk00000003_sig000002c1 : STD_LOGIC; 
  signal blk00000003_sig000002c0 : STD_LOGIC; 
  signal blk00000003_sig000002bf : STD_LOGIC; 
  signal blk00000003_sig000002be : STD_LOGIC; 
  signal blk00000003_sig000002bd : STD_LOGIC; 
  signal blk00000003_sig000002bc : STD_LOGIC; 
  signal blk00000003_sig000002bb : STD_LOGIC; 
  signal blk00000003_sig000002ba : STD_LOGIC; 
  signal blk00000003_sig000002b9 : STD_LOGIC; 
  signal blk00000003_sig000002b8 : STD_LOGIC; 
  signal blk00000003_sig000002b7 : STD_LOGIC; 
  signal blk00000003_sig000002b6 : STD_LOGIC; 
  signal blk00000003_sig000002b5 : STD_LOGIC; 
  signal blk00000003_sig000002b4 : STD_LOGIC; 
  signal blk00000003_sig000002b3 : STD_LOGIC; 
  signal blk00000003_sig000002b2 : STD_LOGIC; 
  signal blk00000003_sig000002b1 : STD_LOGIC; 
  signal blk00000003_sig000002b0 : STD_LOGIC; 
  signal blk00000003_sig000002af : STD_LOGIC; 
  signal blk00000003_sig000002ae : STD_LOGIC; 
  signal blk00000003_sig000002ad : STD_LOGIC; 
  signal blk00000003_sig000002ac : STD_LOGIC; 
  signal blk00000003_sig000002ab : STD_LOGIC; 
  signal blk00000003_sig000002aa : STD_LOGIC; 
  signal blk00000003_sig000002a9 : STD_LOGIC; 
  signal blk00000003_sig000002a8 : STD_LOGIC; 
  signal blk00000003_sig000002a7 : STD_LOGIC; 
  signal blk00000003_sig000002a6 : STD_LOGIC; 
  signal blk00000003_sig000002a5 : STD_LOGIC; 
  signal blk00000003_sig000002a4 : STD_LOGIC; 
  signal blk00000003_sig000002a3 : STD_LOGIC; 
  signal blk00000003_sig000002a2 : STD_LOGIC; 
  signal blk00000003_sig000002a1 : STD_LOGIC; 
  signal blk00000003_sig000002a0 : STD_LOGIC; 
  signal blk00000003_sig0000029f : STD_LOGIC; 
  signal blk00000003_sig0000029e : STD_LOGIC; 
  signal blk00000003_sig0000029d : STD_LOGIC; 
  signal blk00000003_sig0000029c : STD_LOGIC; 
  signal blk00000003_sig0000029b : STD_LOGIC; 
  signal blk00000003_sig0000029a : STD_LOGIC; 
  signal blk00000003_sig00000299 : STD_LOGIC; 
  signal blk00000003_sig00000298 : STD_LOGIC; 
  signal blk00000003_sig00000297 : STD_LOGIC; 
  signal blk00000003_sig00000296 : STD_LOGIC; 
  signal blk00000003_sig00000295 : STD_LOGIC; 
  signal blk00000003_sig00000294 : STD_LOGIC; 
  signal blk00000003_sig00000293 : STD_LOGIC; 
  signal blk00000003_sig00000292 : STD_LOGIC; 
  signal blk00000003_sig00000291 : STD_LOGIC; 
  signal blk00000003_sig00000290 : STD_LOGIC; 
  signal blk00000003_sig0000028f : STD_LOGIC; 
  signal blk00000003_sig0000028e : STD_LOGIC; 
  signal blk00000003_sig0000028d : STD_LOGIC; 
  signal blk00000003_sig0000028c : STD_LOGIC; 
  signal blk00000003_sig0000028b : STD_LOGIC; 
  signal blk00000003_sig0000028a : STD_LOGIC; 
  signal blk00000003_sig00000289 : STD_LOGIC; 
  signal blk00000003_sig00000288 : STD_LOGIC; 
  signal blk00000003_sig00000287 : STD_LOGIC; 
  signal blk00000003_sig00000286 : STD_LOGIC; 
  signal blk00000003_sig00000285 : STD_LOGIC; 
  signal blk00000003_sig00000284 : STD_LOGIC; 
  signal blk00000003_sig00000283 : STD_LOGIC; 
  signal blk00000003_sig00000282 : STD_LOGIC; 
  signal blk00000003_sig00000281 : STD_LOGIC; 
  signal blk00000003_sig00000280 : STD_LOGIC; 
  signal blk00000003_sig0000027f : STD_LOGIC; 
  signal blk00000003_sig0000027e : STD_LOGIC; 
  signal blk00000003_sig0000027d : STD_LOGIC; 
  signal blk00000003_sig0000027c : STD_LOGIC; 
  signal blk00000003_sig0000027b : STD_LOGIC; 
  signal blk00000003_sig0000027a : STD_LOGIC; 
  signal blk00000003_sig00000279 : STD_LOGIC; 
  signal blk00000003_sig00000278 : STD_LOGIC; 
  signal blk00000003_sig00000277 : STD_LOGIC; 
  signal blk00000003_sig00000276 : STD_LOGIC; 
  signal blk00000003_sig00000275 : STD_LOGIC; 
  signal blk00000003_sig00000274 : STD_LOGIC; 
  signal blk00000003_sig00000273 : STD_LOGIC; 
  signal blk00000003_sig00000272 : STD_LOGIC; 
  signal blk00000003_sig00000271 : STD_LOGIC; 
  signal blk00000003_sig00000270 : STD_LOGIC; 
  signal blk00000003_sig0000026f : STD_LOGIC; 
  signal blk00000003_sig0000026e : STD_LOGIC; 
  signal blk00000003_sig0000026d : STD_LOGIC; 
  signal blk00000003_sig0000026c : STD_LOGIC; 
  signal blk00000003_sig0000026b : STD_LOGIC; 
  signal blk00000003_sig0000026a : STD_LOGIC; 
  signal blk00000003_sig00000269 : STD_LOGIC; 
  signal blk00000003_sig00000268 : STD_LOGIC; 
  signal blk00000003_sig00000267 : STD_LOGIC; 
  signal blk00000003_sig00000266 : STD_LOGIC; 
  signal blk00000003_sig00000265 : STD_LOGIC; 
  signal blk00000003_sig00000264 : STD_LOGIC; 
  signal blk00000003_sig00000263 : STD_LOGIC; 
  signal blk00000003_sig00000262 : STD_LOGIC; 
  signal blk00000003_sig00000261 : STD_LOGIC; 
  signal blk00000003_sig00000260 : STD_LOGIC; 
  signal blk00000003_sig0000025f : STD_LOGIC; 
  signal blk00000003_sig0000025e : STD_LOGIC; 
  signal blk00000003_sig0000025d : STD_LOGIC; 
  signal blk00000003_sig0000025c : STD_LOGIC; 
  signal blk00000003_sig0000025b : STD_LOGIC; 
  signal blk00000003_sig0000025a : STD_LOGIC; 
  signal blk00000003_sig00000259 : STD_LOGIC; 
  signal blk00000003_sig00000258 : STD_LOGIC; 
  signal blk00000003_sig00000257 : STD_LOGIC; 
  signal blk00000003_sig00000256 : STD_LOGIC; 
  signal blk00000003_sig00000255 : STD_LOGIC; 
  signal blk00000003_sig00000254 : STD_LOGIC; 
  signal blk00000003_sig00000253 : STD_LOGIC; 
  signal blk00000003_sig00000252 : STD_LOGIC; 
  signal blk00000003_sig00000251 : STD_LOGIC; 
  signal blk00000003_sig00000250 : STD_LOGIC; 
  signal blk00000003_sig0000024f : STD_LOGIC; 
  signal blk00000003_sig0000024e : STD_LOGIC; 
  signal blk00000003_sig0000024d : STD_LOGIC; 
  signal blk00000003_sig0000024c : STD_LOGIC; 
  signal blk00000003_sig0000024b : STD_LOGIC; 
  signal blk00000003_sig0000024a : STD_LOGIC; 
  signal blk00000003_sig00000249 : STD_LOGIC; 
  signal blk00000003_sig00000248 : STD_LOGIC; 
  signal blk00000003_sig00000247 : STD_LOGIC; 
  signal blk00000003_sig00000246 : STD_LOGIC; 
  signal blk00000003_sig00000245 : STD_LOGIC; 
  signal blk00000003_sig00000244 : STD_LOGIC; 
  signal blk00000003_sig00000243 : STD_LOGIC; 
  signal blk00000003_sig00000242 : STD_LOGIC; 
  signal blk00000003_sig00000241 : STD_LOGIC; 
  signal blk00000003_sig00000240 : STD_LOGIC; 
  signal blk00000003_sig0000023f : STD_LOGIC; 
  signal blk00000003_sig0000023e : STD_LOGIC; 
  signal blk00000003_sig0000023d : STD_LOGIC; 
  signal blk00000003_sig0000023c : STD_LOGIC; 
  signal blk00000003_sig0000023b : STD_LOGIC; 
  signal blk00000003_sig0000023a : STD_LOGIC; 
  signal blk00000003_sig00000239 : STD_LOGIC; 
  signal blk00000003_sig00000238 : STD_LOGIC; 
  signal blk00000003_sig00000237 : STD_LOGIC; 
  signal blk00000003_sig00000236 : STD_LOGIC; 
  signal blk00000003_sig00000235 : STD_LOGIC; 
  signal blk00000003_sig00000234 : STD_LOGIC; 
  signal blk00000003_sig00000233 : STD_LOGIC; 
  signal blk00000003_sig00000232 : STD_LOGIC; 
  signal blk00000003_sig00000231 : STD_LOGIC; 
  signal blk00000003_sig00000230 : STD_LOGIC; 
  signal blk00000003_sig0000022f : STD_LOGIC; 
  signal blk00000003_sig0000022e : STD_LOGIC; 
  signal blk00000003_sig0000022d : STD_LOGIC; 
  signal blk00000003_sig0000022c : STD_LOGIC; 
  signal blk00000003_sig0000022b : STD_LOGIC; 
  signal blk00000003_sig0000022a : STD_LOGIC; 
  signal blk00000003_sig00000229 : STD_LOGIC; 
  signal blk00000003_sig00000228 : STD_LOGIC; 
  signal blk00000003_sig00000227 : STD_LOGIC; 
  signal blk00000003_sig00000226 : STD_LOGIC; 
  signal blk00000003_sig00000225 : STD_LOGIC; 
  signal blk00000003_sig00000224 : STD_LOGIC; 
  signal blk00000003_sig00000223 : STD_LOGIC; 
  signal blk00000003_sig00000222 : STD_LOGIC; 
  signal blk00000003_sig00000221 : STD_LOGIC; 
  signal blk00000003_sig00000220 : STD_LOGIC; 
  signal blk00000003_sig0000021f : STD_LOGIC; 
  signal blk00000003_sig0000021e : STD_LOGIC; 
  signal blk00000003_sig0000021d : STD_LOGIC; 
  signal blk00000003_sig0000021c : STD_LOGIC; 
  signal blk00000003_sig0000021b : STD_LOGIC; 
  signal blk00000003_sig0000021a : STD_LOGIC; 
  signal blk00000003_sig00000219 : STD_LOGIC; 
  signal blk00000003_sig00000218 : STD_LOGIC; 
  signal blk00000003_sig00000217 : STD_LOGIC; 
  signal blk00000003_sig00000216 : STD_LOGIC; 
  signal blk00000003_sig00000215 : STD_LOGIC; 
  signal blk00000003_sig00000214 : STD_LOGIC; 
  signal blk00000003_sig00000213 : STD_LOGIC; 
  signal blk00000003_sig00000212 : STD_LOGIC; 
  signal blk00000003_sig00000211 : STD_LOGIC; 
  signal blk00000003_sig00000210 : STD_LOGIC; 
  signal blk00000003_sig0000020f : STD_LOGIC; 
  signal blk00000003_sig0000020e : STD_LOGIC; 
  signal blk00000003_sig0000020d : STD_LOGIC; 
  signal blk00000003_sig0000020c : STD_LOGIC; 
  signal blk00000003_sig0000020b : STD_LOGIC; 
  signal blk00000003_sig0000020a : STD_LOGIC; 
  signal blk00000003_sig00000209 : STD_LOGIC; 
  signal blk00000003_sig00000208 : STD_LOGIC; 
  signal blk00000003_sig00000207 : STD_LOGIC; 
  signal blk00000003_sig00000206 : STD_LOGIC; 
  signal blk00000003_sig00000205 : STD_LOGIC; 
  signal blk00000003_sig00000204 : STD_LOGIC; 
  signal blk00000003_sig00000203 : STD_LOGIC; 
  signal blk00000003_sig00000202 : STD_LOGIC; 
  signal blk00000003_sig00000201 : STD_LOGIC; 
  signal blk00000003_sig00000200 : STD_LOGIC; 
  signal blk00000003_sig000001ff : STD_LOGIC; 
  signal blk00000003_sig000001fe : STD_LOGIC; 
  signal blk00000003_sig000001fd : STD_LOGIC; 
  signal blk00000003_sig000001fc : STD_LOGIC; 
  signal blk00000003_sig000001fb : STD_LOGIC; 
  signal blk00000003_sig000001fa : STD_LOGIC; 
  signal blk00000003_sig000001f9 : STD_LOGIC; 
  signal blk00000003_sig000001f8 : STD_LOGIC; 
  signal blk00000003_sig000001f7 : STD_LOGIC; 
  signal blk00000003_sig000001f6 : STD_LOGIC; 
  signal blk00000003_sig000001f5 : STD_LOGIC; 
  signal blk00000003_sig000001f4 : STD_LOGIC; 
  signal blk00000003_sig000001f3 : STD_LOGIC; 
  signal blk00000003_sig000001f2 : STD_LOGIC; 
  signal blk00000003_sig000001f1 : STD_LOGIC; 
  signal blk00000003_sig000001f0 : STD_LOGIC; 
  signal blk00000003_sig000001ef : STD_LOGIC; 
  signal blk00000003_sig000001ee : STD_LOGIC; 
  signal blk00000003_sig000001ed : STD_LOGIC; 
  signal blk00000003_sig000001ec : STD_LOGIC; 
  signal blk00000003_sig000001eb : STD_LOGIC; 
  signal blk00000003_sig000001ea : STD_LOGIC; 
  signal blk00000003_sig000001e9 : STD_LOGIC; 
  signal blk00000003_sig000001e8 : STD_LOGIC; 
  signal blk00000003_sig000001e7 : STD_LOGIC; 
  signal blk00000003_sig000001e6 : STD_LOGIC; 
  signal blk00000003_sig000001e5 : STD_LOGIC; 
  signal blk00000003_sig000001e4 : STD_LOGIC; 
  signal blk00000003_sig000001e3 : STD_LOGIC; 
  signal blk00000003_sig000001e2 : STD_LOGIC; 
  signal blk00000003_sig000001e1 : STD_LOGIC; 
  signal blk00000003_sig000001e0 : STD_LOGIC; 
  signal blk00000003_sig000001df : STD_LOGIC; 
  signal blk00000003_sig000001de : STD_LOGIC; 
  signal blk00000003_sig000001dd : STD_LOGIC; 
  signal blk00000003_sig000001dc : STD_LOGIC; 
  signal blk00000003_sig000001db : STD_LOGIC; 
  signal blk00000003_sig000001da : STD_LOGIC; 
  signal blk00000003_sig000001d9 : STD_LOGIC; 
  signal blk00000003_sig000001d8 : STD_LOGIC; 
  signal blk00000003_sig000001d7 : STD_LOGIC; 
  signal blk00000003_sig000001d6 : STD_LOGIC; 
  signal blk00000003_sig000001d5 : STD_LOGIC; 
  signal blk00000003_sig000001d4 : STD_LOGIC; 
  signal blk00000003_sig000001d3 : STD_LOGIC; 
  signal blk00000003_sig000001d2 : STD_LOGIC; 
  signal blk00000003_sig000001d1 : STD_LOGIC; 
  signal blk00000003_sig000001d0 : STD_LOGIC; 
  signal blk00000003_sig000001cf : STD_LOGIC; 
  signal blk00000003_sig000001ce : STD_LOGIC; 
  signal blk00000003_sig000001cd : STD_LOGIC; 
  signal blk00000003_sig000001cc : STD_LOGIC; 
  signal blk00000003_sig000001cb : STD_LOGIC; 
  signal blk00000003_sig000001ca : STD_LOGIC; 
  signal blk00000003_sig000001c9 : STD_LOGIC; 
  signal blk00000003_sig000001c8 : STD_LOGIC; 
  signal blk00000003_sig000001c7 : STD_LOGIC; 
  signal blk00000003_sig000001c6 : STD_LOGIC; 
  signal blk00000003_sig000001c5 : STD_LOGIC; 
  signal blk00000003_sig000001c4 : STD_LOGIC; 
  signal blk00000003_sig000001c3 : STD_LOGIC; 
  signal blk00000003_sig000001c2 : STD_LOGIC; 
  signal blk00000003_sig000001c1 : STD_LOGIC; 
  signal blk00000003_sig000001c0 : STD_LOGIC; 
  signal blk00000003_sig000001bf : STD_LOGIC; 
  signal blk00000003_sig000001be : STD_LOGIC; 
  signal blk00000003_sig000001bd : STD_LOGIC; 
  signal blk00000003_sig000001bc : STD_LOGIC; 
  signal blk00000003_sig000001bb : STD_LOGIC; 
  signal blk00000003_sig000001ba : STD_LOGIC; 
  signal blk00000003_sig000001b9 : STD_LOGIC; 
  signal blk00000003_sig000001b8 : STD_LOGIC; 
  signal blk00000003_sig000001b7 : STD_LOGIC; 
  signal blk00000003_sig000001b6 : STD_LOGIC; 
  signal blk00000003_sig000001b5 : STD_LOGIC; 
  signal blk00000003_sig000001b4 : STD_LOGIC; 
  signal blk00000003_sig000001b3 : STD_LOGIC; 
  signal blk00000003_sig000001b2 : STD_LOGIC; 
  signal blk00000003_sig000001b1 : STD_LOGIC; 
  signal blk00000003_sig000001b0 : STD_LOGIC; 
  signal blk00000003_sig000001af : STD_LOGIC; 
  signal blk00000003_sig000001ae : STD_LOGIC; 
  signal blk00000003_sig000001ad : STD_LOGIC; 
  signal blk00000003_sig000001ac : STD_LOGIC; 
  signal blk00000003_sig000001ab : STD_LOGIC; 
  signal blk00000003_sig000001aa : STD_LOGIC; 
  signal blk00000003_sig000001a9 : STD_LOGIC; 
  signal blk00000003_sig000001a8 : STD_LOGIC; 
  signal blk00000003_sig000001a7 : STD_LOGIC; 
  signal blk00000003_sig000001a6 : STD_LOGIC; 
  signal blk00000003_sig000001a5 : STD_LOGIC; 
  signal blk00000003_sig000001a4 : STD_LOGIC; 
  signal blk00000003_sig000001a3 : STD_LOGIC; 
  signal blk00000003_sig000001a2 : STD_LOGIC; 
  signal blk00000003_sig000001a1 : STD_LOGIC; 
  signal blk00000003_sig000001a0 : STD_LOGIC; 
  signal blk00000003_sig0000019f : STD_LOGIC; 
  signal blk00000003_sig0000019e : STD_LOGIC; 
  signal blk00000003_sig0000019d : STD_LOGIC; 
  signal blk00000003_sig0000019c : STD_LOGIC; 
  signal blk00000003_sig0000019b : STD_LOGIC; 
  signal blk00000003_sig0000019a : STD_LOGIC; 
  signal blk00000003_sig00000199 : STD_LOGIC; 
  signal blk00000003_sig00000198 : STD_LOGIC; 
  signal blk00000003_sig00000197 : STD_LOGIC; 
  signal blk00000003_sig00000196 : STD_LOGIC; 
  signal blk00000003_sig00000195 : STD_LOGIC; 
  signal blk00000003_sig00000194 : STD_LOGIC; 
  signal blk00000003_sig00000193 : STD_LOGIC; 
  signal blk00000003_sig00000192 : STD_LOGIC; 
  signal blk00000003_sig00000191 : STD_LOGIC; 
  signal blk00000003_sig00000190 : STD_LOGIC; 
  signal blk00000003_sig0000018f : STD_LOGIC; 
  signal blk00000003_sig0000018e : STD_LOGIC; 
  signal blk00000003_sig0000018d : STD_LOGIC; 
  signal blk00000003_sig0000018c : STD_LOGIC; 
  signal blk00000003_sig0000018b : STD_LOGIC; 
  signal blk00000003_sig0000018a : STD_LOGIC; 
  signal blk00000003_sig00000189 : STD_LOGIC; 
  signal blk00000003_sig00000188 : STD_LOGIC; 
  signal blk00000003_sig00000187 : STD_LOGIC; 
  signal blk00000003_sig00000186 : STD_LOGIC; 
  signal blk00000003_sig00000185 : STD_LOGIC; 
  signal blk00000003_sig00000184 : STD_LOGIC; 
  signal blk00000003_sig00000183 : STD_LOGIC; 
  signal blk00000003_sig00000182 : STD_LOGIC; 
  signal blk00000003_sig00000181 : STD_LOGIC; 
  signal blk00000003_sig00000180 : STD_LOGIC; 
  signal blk00000003_sig0000017f : STD_LOGIC; 
  signal blk00000003_sig0000017e : STD_LOGIC; 
  signal blk00000003_sig0000017d : STD_LOGIC; 
  signal blk00000003_sig0000017c : STD_LOGIC; 
  signal blk00000003_sig0000017b : STD_LOGIC; 
  signal blk00000003_sig0000017a : STD_LOGIC; 
  signal blk00000003_sig00000179 : STD_LOGIC; 
  signal blk00000003_sig00000178 : STD_LOGIC; 
  signal blk00000003_sig00000177 : STD_LOGIC; 
  signal blk00000003_sig00000176 : STD_LOGIC; 
  signal blk00000003_sig00000175 : STD_LOGIC; 
  signal blk00000003_sig00000174 : STD_LOGIC; 
  signal blk00000003_sig00000173 : STD_LOGIC; 
  signal blk00000003_sig00000172 : STD_LOGIC; 
  signal blk00000003_sig00000171 : STD_LOGIC; 
  signal blk00000003_sig00000170 : STD_LOGIC; 
  signal blk00000003_sig0000016f : STD_LOGIC; 
  signal blk00000003_sig0000016e : STD_LOGIC; 
  signal blk00000003_sig0000016d : STD_LOGIC; 
  signal blk00000003_sig0000016c : STD_LOGIC; 
  signal blk00000003_sig0000016b : STD_LOGIC; 
  signal blk00000003_sig0000016a : STD_LOGIC; 
  signal blk00000003_sig00000169 : STD_LOGIC; 
  signal blk00000003_sig00000168 : STD_LOGIC; 
  signal blk00000003_sig00000167 : STD_LOGIC; 
  signal blk00000003_sig00000166 : STD_LOGIC; 
  signal blk00000003_sig00000165 : STD_LOGIC; 
  signal blk00000003_sig00000164 : STD_LOGIC; 
  signal blk00000003_sig00000163 : STD_LOGIC; 
  signal blk00000003_sig00000162 : STD_LOGIC; 
  signal blk00000003_sig00000161 : STD_LOGIC; 
  signal blk00000003_sig00000160 : STD_LOGIC; 
  signal blk00000003_sig0000015f : STD_LOGIC; 
  signal blk00000003_sig0000015e : STD_LOGIC; 
  signal blk00000003_sig0000015d : STD_LOGIC; 
  signal blk00000003_sig0000015c : STD_LOGIC; 
  signal blk00000003_sig0000015b : STD_LOGIC; 
  signal blk00000003_sig0000015a : STD_LOGIC; 
  signal blk00000003_sig00000159 : STD_LOGIC; 
  signal blk00000003_sig00000158 : STD_LOGIC; 
  signal blk00000003_sig00000157 : STD_LOGIC; 
  signal blk00000003_sig00000156 : STD_LOGIC; 
  signal blk00000003_sig00000155 : STD_LOGIC; 
  signal blk00000003_sig00000154 : STD_LOGIC; 
  signal blk00000003_sig00000153 : STD_LOGIC; 
  signal blk00000003_sig00000152 : STD_LOGIC; 
  signal blk00000003_sig00000151 : STD_LOGIC; 
  signal blk00000003_sig00000150 : STD_LOGIC; 
  signal blk00000003_sig0000014f : STD_LOGIC; 
  signal blk00000003_sig0000014e : STD_LOGIC; 
  signal blk00000003_sig0000014d : STD_LOGIC; 
  signal blk00000003_sig0000014c : STD_LOGIC; 
  signal blk00000003_sig0000014b : STD_LOGIC; 
  signal blk00000003_sig0000014a : STD_LOGIC; 
  signal blk00000003_sig00000149 : STD_LOGIC; 
  signal blk00000003_sig00000148 : STD_LOGIC; 
  signal blk00000003_sig00000147 : STD_LOGIC; 
  signal blk00000003_sig00000146 : STD_LOGIC; 
  signal blk00000003_sig00000145 : STD_LOGIC; 
  signal blk00000003_sig00000144 : STD_LOGIC; 
  signal blk00000003_sig00000143 : STD_LOGIC; 
  signal blk00000003_sig00000142 : STD_LOGIC; 
  signal blk00000003_sig00000141 : STD_LOGIC; 
  signal blk00000003_sig00000140 : STD_LOGIC; 
  signal blk00000003_sig0000013f : STD_LOGIC; 
  signal blk00000003_sig0000013e : STD_LOGIC; 
  signal blk00000003_sig0000013d : STD_LOGIC; 
  signal blk00000003_sig0000013c : STD_LOGIC; 
  signal blk00000003_sig0000013b : STD_LOGIC; 
  signal blk00000003_sig0000013a : STD_LOGIC; 
  signal blk00000003_sig00000139 : STD_LOGIC; 
  signal blk00000003_sig00000138 : STD_LOGIC; 
  signal blk00000003_sig00000137 : STD_LOGIC; 
  signal blk00000003_sig00000136 : STD_LOGIC; 
  signal blk00000003_sig00000135 : STD_LOGIC; 
  signal blk00000003_sig00000134 : STD_LOGIC; 
  signal blk00000003_sig00000133 : STD_LOGIC; 
  signal blk00000003_sig00000132 : STD_LOGIC; 
  signal blk00000003_sig00000131 : STD_LOGIC; 
  signal blk00000003_sig00000130 : STD_LOGIC; 
  signal blk00000003_sig0000012f : STD_LOGIC; 
  signal blk00000003_sig0000012e : STD_LOGIC; 
  signal blk00000003_sig0000012d : STD_LOGIC; 
  signal blk00000003_sig0000012c : STD_LOGIC; 
  signal blk00000003_sig0000012b : STD_LOGIC; 
  signal blk00000003_sig0000012a : STD_LOGIC; 
  signal blk00000003_sig00000129 : STD_LOGIC; 
  signal blk00000003_sig00000128 : STD_LOGIC; 
  signal blk00000003_sig00000127 : STD_LOGIC; 
  signal blk00000003_sig00000126 : STD_LOGIC; 
  signal blk00000003_sig00000125 : STD_LOGIC; 
  signal blk00000003_sig00000124 : STD_LOGIC; 
  signal blk00000003_sig00000123 : STD_LOGIC; 
  signal blk00000003_sig00000122 : STD_LOGIC; 
  signal blk00000003_sig00000121 : STD_LOGIC; 
  signal blk00000003_sig00000120 : STD_LOGIC; 
  signal blk00000003_sig0000011f : STD_LOGIC; 
  signal blk00000003_sig0000011e : STD_LOGIC; 
  signal blk00000003_sig0000011d : STD_LOGIC; 
  signal blk00000003_sig0000011c : STD_LOGIC; 
  signal blk00000003_sig0000011b : STD_LOGIC; 
  signal blk00000003_sig0000011a : STD_LOGIC; 
  signal blk00000003_sig00000119 : STD_LOGIC; 
  signal blk00000003_sig00000118 : STD_LOGIC; 
  signal blk00000003_sig00000117 : STD_LOGIC; 
  signal blk00000003_sig00000116 : STD_LOGIC; 
  signal blk00000003_sig00000115 : STD_LOGIC; 
  signal blk00000003_sig00000114 : STD_LOGIC; 
  signal blk00000003_sig00000113 : STD_LOGIC; 
  signal blk00000003_sig00000112 : STD_LOGIC; 
  signal blk00000003_sig00000111 : STD_LOGIC; 
  signal blk00000003_sig00000110 : STD_LOGIC; 
  signal blk00000003_sig0000010f : STD_LOGIC; 
  signal blk00000003_sig0000010e : STD_LOGIC; 
  signal blk00000003_sig0000010d : STD_LOGIC; 
  signal blk00000003_sig0000010c : STD_LOGIC; 
  signal blk00000003_sig0000010b : STD_LOGIC; 
  signal blk00000003_sig0000010a : STD_LOGIC; 
  signal blk00000003_sig00000109 : STD_LOGIC; 
  signal blk00000003_sig00000108 : STD_LOGIC; 
  signal blk00000003_sig00000107 : STD_LOGIC; 
  signal blk00000003_sig00000106 : STD_LOGIC; 
  signal blk00000003_sig00000105 : STD_LOGIC; 
  signal blk00000003_sig00000104 : STD_LOGIC; 
  signal blk00000003_sig00000103 : STD_LOGIC; 
  signal blk00000003_sig00000102 : STD_LOGIC; 
  signal blk00000003_sig00000101 : STD_LOGIC; 
  signal blk00000003_sig00000100 : STD_LOGIC; 
  signal blk00000003_sig000000ff : STD_LOGIC; 
  signal blk00000003_sig000000fe : STD_LOGIC; 
  signal blk00000003_sig000000fd : STD_LOGIC; 
  signal blk00000003_sig000000fc : STD_LOGIC; 
  signal blk00000003_sig000000fb : STD_LOGIC; 
  signal blk00000003_sig000000fa : STD_LOGIC; 
  signal blk00000003_sig000000f9 : STD_LOGIC; 
  signal blk00000003_sig000000f8 : STD_LOGIC; 
  signal blk00000003_sig000000f7 : STD_LOGIC; 
  signal blk00000003_sig000000f6 : STD_LOGIC; 
  signal blk00000003_sig000000f5 : STD_LOGIC; 
  signal blk00000003_sig000000f4 : STD_LOGIC; 
  signal blk00000003_sig000000f3 : STD_LOGIC; 
  signal blk00000003_sig000000f2 : STD_LOGIC; 
  signal blk00000003_sig000000f1 : STD_LOGIC; 
  signal blk00000003_sig000000f0 : STD_LOGIC; 
  signal blk00000003_sig000000ef : STD_LOGIC; 
  signal blk00000003_sig000000ee : STD_LOGIC; 
  signal blk00000003_sig000000ed : STD_LOGIC; 
  signal blk00000003_sig000000ec : STD_LOGIC; 
  signal blk00000003_sig000000eb : STD_LOGIC; 
  signal blk00000003_sig000000ea : STD_LOGIC; 
  signal blk00000003_sig000000e9 : STD_LOGIC; 
  signal blk00000003_sig000000e8 : STD_LOGIC; 
  signal blk00000003_sig000000e7 : STD_LOGIC; 
  signal blk00000003_sig000000e6 : STD_LOGIC; 
  signal blk00000003_sig000000e5 : STD_LOGIC; 
  signal blk00000003_sig000000e4 : STD_LOGIC; 
  signal blk00000003_sig000000e3 : STD_LOGIC; 
  signal blk00000003_sig000000e2 : STD_LOGIC; 
  signal blk00000003_sig000000e1 : STD_LOGIC; 
  signal blk00000003_sig000000e0 : STD_LOGIC; 
  signal blk00000003_sig000000df : STD_LOGIC; 
  signal blk00000003_sig000000de : STD_LOGIC; 
  signal blk00000003_sig000000dd : STD_LOGIC; 
  signal blk00000003_sig000000dc : STD_LOGIC; 
  signal blk00000003_sig000000db : STD_LOGIC; 
  signal blk00000003_sig000000da : STD_LOGIC; 
  signal blk00000003_sig000000d9 : STD_LOGIC; 
  signal blk00000003_sig000000d8 : STD_LOGIC; 
  signal blk00000003_sig000000d7 : STD_LOGIC; 
  signal blk00000003_sig000000d6 : STD_LOGIC; 
  signal blk00000003_sig000000d5 : STD_LOGIC; 
  signal blk00000003_sig000000d4 : STD_LOGIC; 
  signal blk00000003_sig000000d3 : STD_LOGIC; 
  signal blk00000003_sig000000d2 : STD_LOGIC; 
  signal blk00000003_sig000000d1 : STD_LOGIC; 
  signal blk00000003_sig000000d0 : STD_LOGIC; 
  signal blk00000003_sig000000cf : STD_LOGIC; 
  signal blk00000003_sig000000ce : STD_LOGIC; 
  signal blk00000003_sig000000cd : STD_LOGIC; 
  signal blk00000003_sig000000cc : STD_LOGIC; 
  signal blk00000003_sig000000cb : STD_LOGIC; 
  signal blk00000003_sig000000ca : STD_LOGIC; 
  signal blk00000003_sig000000c9 : STD_LOGIC; 
  signal blk00000003_sig000000c8 : STD_LOGIC; 
  signal blk00000003_sig000000c7 : STD_LOGIC; 
  signal blk00000003_sig000000c6 : STD_LOGIC; 
  signal blk00000003_sig000000c5 : STD_LOGIC; 
  signal blk00000003_sig000000c4 : STD_LOGIC; 
  signal blk00000003_sig000000c3 : STD_LOGIC; 
  signal blk00000003_sig000000c2 : STD_LOGIC; 
  signal blk00000003_sig000000c1 : STD_LOGIC; 
  signal blk00000003_sig000000c0 : STD_LOGIC; 
  signal blk00000003_sig000000bf : STD_LOGIC; 
  signal blk00000003_sig000000be : STD_LOGIC; 
  signal blk00000003_sig000000bd : STD_LOGIC; 
  signal blk00000003_sig000000bc : STD_LOGIC; 
  signal blk00000003_sig000000bb : STD_LOGIC; 
  signal blk00000003_sig000000ba : STD_LOGIC; 
  signal blk00000003_sig000000b9 : STD_LOGIC; 
  signal blk00000003_sig000000b8 : STD_LOGIC; 
  signal blk00000003_sig000000b7 : STD_LOGIC; 
  signal blk00000003_sig000000b6 : STD_LOGIC; 
  signal blk00000003_sig000000b5 : STD_LOGIC; 
  signal blk00000003_sig000000b4 : STD_LOGIC; 
  signal blk00000003_sig000000b3 : STD_LOGIC; 
  signal blk00000003_sig000000b2 : STD_LOGIC; 
  signal blk00000003_sig000000b1 : STD_LOGIC; 
  signal blk00000003_sig000000b0 : STD_LOGIC; 
  signal blk00000003_sig000000af : STD_LOGIC; 
  signal blk00000003_sig000000ae : STD_LOGIC; 
  signal blk00000003_sig000000ad : STD_LOGIC; 
  signal blk00000003_sig000000ac : STD_LOGIC; 
  signal blk00000003_sig000000ab : STD_LOGIC; 
  signal blk00000003_sig000000aa : STD_LOGIC; 
  signal blk00000003_sig000000a9 : STD_LOGIC; 
  signal blk00000003_sig000000a8 : STD_LOGIC; 
  signal blk00000003_sig000000a7 : STD_LOGIC; 
  signal blk00000003_sig000000a6 : STD_LOGIC; 
  signal blk00000003_sig000000a5 : STD_LOGIC; 
  signal blk00000003_sig000000a4 : STD_LOGIC; 
  signal blk00000003_sig000000a3 : STD_LOGIC; 
  signal blk00000003_sig000000a2 : STD_LOGIC; 
  signal blk00000003_sig000000a1 : STD_LOGIC; 
  signal blk00000003_sig000000a0 : STD_LOGIC; 
  signal blk00000003_sig0000009f : STD_LOGIC; 
  signal blk00000003_sig0000009e : STD_LOGIC; 
  signal blk00000003_sig0000009d : STD_LOGIC; 
  signal blk00000003_sig0000009c : STD_LOGIC; 
  signal blk00000003_sig0000009b : STD_LOGIC; 
  signal blk00000003_sig0000009a : STD_LOGIC; 
  signal blk00000003_sig00000099 : STD_LOGIC; 
  signal blk00000003_sig00000098 : STD_LOGIC; 
  signal blk00000003_sig00000097 : STD_LOGIC; 
  signal blk00000003_sig00000096 : STD_LOGIC; 
  signal blk00000003_sig00000095 : STD_LOGIC; 
  signal blk00000003_sig00000094 : STD_LOGIC; 
  signal blk00000003_sig00000093 : STD_LOGIC; 
  signal blk00000003_sig00000092 : STD_LOGIC; 
  signal blk00000003_sig00000091 : STD_LOGIC; 
  signal blk00000003_sig00000090 : STD_LOGIC; 
  signal blk00000003_sig0000008f : STD_LOGIC; 
  signal blk00000003_sig0000008e : STD_LOGIC; 
  signal blk00000003_sig0000008d : STD_LOGIC; 
  signal blk00000003_sig0000008c : STD_LOGIC; 
  signal blk00000003_sig0000008b : STD_LOGIC; 
  signal blk00000003_sig0000008a : STD_LOGIC; 
  signal blk00000003_sig00000089 : STD_LOGIC; 
  signal blk00000003_sig00000088 : STD_LOGIC; 
  signal blk00000003_sig00000087 : STD_LOGIC; 
  signal blk00000003_sig00000086 : STD_LOGIC; 
  signal blk00000003_sig00000085 : STD_LOGIC; 
  signal blk00000003_sig00000084 : STD_LOGIC; 
  signal blk00000003_sig00000083 : STD_LOGIC; 
  signal blk00000003_sig00000082 : STD_LOGIC; 
  signal blk00000003_sig00000081 : STD_LOGIC; 
  signal blk00000003_sig00000080 : STD_LOGIC; 
  signal blk00000003_sig0000007f : STD_LOGIC; 
  signal blk00000003_sig0000007e : STD_LOGIC; 
  signal blk00000003_sig0000007d : STD_LOGIC; 
  signal blk00000003_sig0000007c : STD_LOGIC; 
  signal blk00000003_sig0000007b : STD_LOGIC; 
  signal blk00000003_sig0000007a : STD_LOGIC; 
  signal blk00000003_sig00000079 : STD_LOGIC; 
  signal blk00000003_sig00000078 : STD_LOGIC; 
  signal blk00000003_sig00000077 : STD_LOGIC; 
  signal blk00000003_sig00000076 : STD_LOGIC; 
  signal blk00000003_sig00000075 : STD_LOGIC; 
  signal blk00000003_sig00000074 : STD_LOGIC; 
  signal blk00000003_sig00000073 : STD_LOGIC; 
  signal blk00000003_sig00000072 : STD_LOGIC; 
  signal blk00000003_sig00000071 : STD_LOGIC; 
  signal blk00000003_sig00000070 : STD_LOGIC; 
  signal blk00000003_sig0000006f : STD_LOGIC; 
  signal blk00000003_sig0000006e : STD_LOGIC; 
  signal blk00000003_sig0000006d : STD_LOGIC; 
  signal blk00000003_sig0000006c : STD_LOGIC; 
  signal blk00000003_sig0000006b : STD_LOGIC; 
  signal blk00000003_sig0000006a : STD_LOGIC; 
  signal blk00000003_sig00000069 : STD_LOGIC; 
  signal blk00000003_sig00000068 : STD_LOGIC; 
  signal blk00000003_sig00000067 : STD_LOGIC; 
  signal blk00000003_sig00000066 : STD_LOGIC; 
  signal blk00000003_sig00000065 : STD_LOGIC; 
  signal blk00000003_sig00000064 : STD_LOGIC; 
  signal blk00000003_sig00000063 : STD_LOGIC; 
  signal blk00000003_sig00000062 : STD_LOGIC; 
  signal blk00000003_sig00000061 : STD_LOGIC; 
  signal blk00000003_sig00000060 : STD_LOGIC; 
  signal blk00000003_sig0000005f : STD_LOGIC; 
  signal blk00000003_sig0000005e : STD_LOGIC; 
  signal blk00000003_sig0000005d : STD_LOGIC; 
  signal blk00000003_sig0000005c : STD_LOGIC; 
  signal blk00000003_sig0000005b : STD_LOGIC; 
  signal blk00000003_sig0000005a : STD_LOGIC; 
  signal blk00000003_sig00000059 : STD_LOGIC; 
  signal blk00000003_sig00000058 : STD_LOGIC; 
  signal blk00000003_sig00000057 : STD_LOGIC; 
  signal blk00000003_sig00000056 : STD_LOGIC; 
  signal blk00000003_sig00000055 : STD_LOGIC; 
  signal blk00000003_sig00000054 : STD_LOGIC; 
  signal blk00000003_sig00000053 : STD_LOGIC; 
  signal blk00000003_sig00000052 : STD_LOGIC; 
  signal blk00000003_sig00000051 : STD_LOGIC; 
  signal blk00000003_sig0000004f : STD_LOGIC; 
  signal NLW_blk00000001_P_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000002_G_UNCONNECTED : STD_LOGIC; 
  signal NLW_blk00000003_blk0000014f_O_UNCONNECTED : STD_LOGIC; 
begin
  rfd <= NlwRenamedSig_OI_rfd;
  blk00000001 : VCC
    port map (
      P => NLW_blk00000001_P_UNCONNECTED
    );
  blk00000002 : GND
    port map (
      G => NLW_blk00000002_G_UNCONNECTED
    );
  blk00000003_blk000008ec : INV
    port map (
      I => blk00000003_sig0000009c,
      O => blk00000003_sig000001a0
    );
  blk00000003_blk000008eb : INV
    port map (
      I => blk00000003_sig0000009b,
      O => blk00000003_sig000001a3
    );
  blk00000003_blk000008ea : INV
    port map (
      I => blk00000003_sig0000009a,
      O => blk00000003_sig000001a6
    );
  blk00000003_blk000008e9 : INV
    port map (
      I => blk00000003_sig00000099,
      O => blk00000003_sig000001a9
    );
  blk00000003_blk000008e8 : INV
    port map (
      I => blk00000003_sig00000098,
      O => blk00000003_sig000001ac
    );
  blk00000003_blk000008e7 : INV
    port map (
      I => blk00000003_sig000008d4,
      O => blk00000003_sig0000015d
    );
  blk00000003_blk000008e6 : INV
    port map (
      I => blk00000003_sig000008d5,
      O => blk00000003_sig0000015e
    );
  blk00000003_blk000008e5 : INV
    port map (
      I => blk00000003_sig000008d6,
      O => blk00000003_sig0000015f
    );
  blk00000003_blk000008e4 : INV
    port map (
      I => blk00000003_sig000008d7,
      O => blk00000003_sig00000160
    );
  blk00000003_blk000008e3 : INV
    port map (
      I => blk00000003_sig000008d8,
      O => blk00000003_sig00000161
    );
  blk00000003_blk000008e2 : INV
    port map (
      I => blk00000003_sig000008d9,
      O => blk00000003_sig00000162
    );
  blk00000003_blk000008e1 : INV
    port map (
      I => blk00000003_sig000008da,
      O => blk00000003_sig00000163
    );
  blk00000003_blk000008e0 : INV
    port map (
      I => blk00000003_sig000008db,
      O => blk00000003_sig00000164
    );
  blk00000003_blk000008df : INV
    port map (
      I => blk00000003_sig000008dc,
      O => blk00000003_sig00000165
    );
  blk00000003_blk000008de : INV
    port map (
      I => blk00000003_sig000008dd,
      O => blk00000003_sig00000166
    );
  blk00000003_blk000008dd : INV
    port map (
      I => blk00000003_sig000008de,
      O => blk00000003_sig00000167
    );
  blk00000003_blk000008dc : INV
    port map (
      I => blk00000003_sig000008df,
      O => blk00000003_sig00000168
    );
  blk00000003_blk000008db : INV
    port map (
      I => blk00000003_sig000008e0,
      O => blk00000003_sig00000169
    );
  blk00000003_blk000008da : INV
    port map (
      I => blk00000003_sig000008e1,
      O => blk00000003_sig0000016a
    );
  blk00000003_blk000008d9 : INV
    port map (
      I => blk00000003_sig000008e2,
      O => blk00000003_sig0000016b
    );
  blk00000003_blk000008d8 : INV
    port map (
      I => blk00000003_sig000008e3,
      O => blk00000003_sig0000016c
    );
  blk00000003_blk000008d7 : INV
    port map (
      I => blk00000003_sig000008e4,
      O => blk00000003_sig0000016d
    );
  blk00000003_blk000008d6 : INV
    port map (
      I => blk00000003_sig000008e5,
      O => blk00000003_sig0000016e
    );
  blk00000003_blk000008d5 : INV
    port map (
      I => blk00000003_sig000008e6,
      O => blk00000003_sig0000016f
    );
  blk00000003_blk000008d4 : INV
    port map (
      I => blk00000003_sig000008e7,
      O => blk00000003_sig00000170
    );
  blk00000003_blk000008d3 : INV
    port map (
      I => blk00000003_sig000008e8,
      O => blk00000003_sig00000171
    );
  blk00000003_blk000008d2 : INV
    port map (
      I => blk00000003_sig000008e9,
      O => blk00000003_sig00000172
    );
  blk00000003_blk000008d1 : INV
    port map (
      I => blk00000003_sig000008ea,
      O => blk00000003_sig00000173
    );
  blk00000003_blk000008d0 : INV
    port map (
      I => blk00000003_sig000008eb,
      O => blk00000003_sig00000174
    );
  blk00000003_blk000008cf : INV
    port map (
      I => blk00000003_sig000008ec,
      O => blk00000003_sig00000175
    );
  blk00000003_blk000008ce : INV
    port map (
      I => blk00000003_sig000008ed,
      O => blk00000003_sig00000176
    );
  blk00000003_blk000008cd : INV
    port map (
      I => blk00000003_sig000008ee,
      O => blk00000003_sig00000177
    );
  blk00000003_blk000008cc : INV
    port map (
      I => blk00000003_sig000008ef,
      O => blk00000003_sig00000178
    );
  blk00000003_blk000008cb : INV
    port map (
      I => blk00000003_sig000008f0,
      O => blk00000003_sig00000179
    );
  blk00000003_blk000008ca : INV
    port map (
      I => blk00000003_sig000008f1,
      O => blk00000003_sig0000017a
    );
  blk00000003_blk000008c9 : INV
    port map (
      I => blk00000003_sig000008f2,
      O => blk00000003_sig0000017b
    );
  blk00000003_blk000008c8 : INV
    port map (
      I => blk00000003_sig0000054a,
      O => blk00000003_sig0000055f
    );
  blk00000003_blk000008c7 : INV
    port map (
      I => blk00000003_sig0000052c,
      O => blk00000003_sig00000541
    );
  blk00000003_blk000008c6 : INV
    port map (
      I => blk00000003_sig0000050e,
      O => blk00000003_sig00000523
    );
  blk00000003_blk000008c5 : INV
    port map (
      I => blk00000003_sig000004f0,
      O => blk00000003_sig00000505
    );
  blk00000003_blk000008c4 : INV
    port map (
      I => blk00000003_sig000004d2,
      O => blk00000003_sig000004e7
    );
  blk00000003_blk000008c3 : INV
    port map (
      I => blk00000003_sig000004b4,
      O => blk00000003_sig000004c9
    );
  blk00000003_blk000008c2 : INV
    port map (
      I => blk00000003_sig00000496,
      O => blk00000003_sig000004ab
    );
  blk00000003_blk000008c1 : INV
    port map (
      I => blk00000003_sig00000477,
      O => blk00000003_sig0000048c
    );
  blk00000003_blk000008c0 : INV
    port map (
      I => blk00000003_sig00000458,
      O => blk00000003_sig0000046d
    );
  blk00000003_blk000008bf : INV
    port map (
      I => blk00000003_sig00000439,
      O => blk00000003_sig0000044e
    );
  blk00000003_blk000008be : INV
    port map (
      I => blk00000003_sig0000041a,
      O => blk00000003_sig0000042f
    );
  blk00000003_blk000008bd : INV
    port map (
      I => blk00000003_sig000003fb,
      O => blk00000003_sig00000410
    );
  blk00000003_blk000008bc : INV
    port map (
      I => blk00000003_sig000003dc,
      O => blk00000003_sig000003f1
    );
  blk00000003_blk000008bb : INV
    port map (
      I => blk00000003_sig000003bd,
      O => blk00000003_sig000003d2
    );
  blk00000003_blk000008ba : INV
    port map (
      I => blk00000003_sig0000039e,
      O => blk00000003_sig000003b3
    );
  blk00000003_blk000008b9 : INV
    port map (
      I => blk00000003_sig0000037f,
      O => blk00000003_sig00000394
    );
  blk00000003_blk000008b8 : INV
    port map (
      I => blk00000003_sig00000360,
      O => blk00000003_sig00000375
    );
  blk00000003_blk000008b7 : INV
    port map (
      I => blk00000003_sig00000341,
      O => blk00000003_sig00000356
    );
  blk00000003_blk000008b6 : INV
    port map (
      I => blk00000003_sig00000322,
      O => blk00000003_sig00000337
    );
  blk00000003_blk000008b5 : INV
    port map (
      I => blk00000003_sig00000303,
      O => blk00000003_sig00000318
    );
  blk00000003_blk000008b4 : INV
    port map (
      I => blk00000003_sig000002e4,
      O => blk00000003_sig000002f9
    );
  blk00000003_blk000008b3 : INV
    port map (
      I => blk00000003_sig000002c5,
      O => blk00000003_sig000002da
    );
  blk00000003_blk000008b2 : INV
    port map (
      I => blk00000003_sig000002a6,
      O => blk00000003_sig000002bb
    );
  blk00000003_blk000008b1 : INV
    port map (
      I => blk00000003_sig00000287,
      O => blk00000003_sig0000029c
    );
  blk00000003_blk000008b0 : INV
    port map (
      I => blk00000003_sig0000008e,
      O => blk00000003_sig0000027d
    );
  blk00000003_blk000008af : INV
    port map (
      I => blk00000003_sig00000073,
      O => blk00000003_sig0000025f
    );
  blk00000003_blk000008ae : INV
    port map (
      I => blk00000003_sig0000007f,
      O => blk00000003_sig00000241
    );
  blk00000003_blk000008ad : INV
    port map (
      I => blk00000003_sig00000084,
      O => blk00000003_sig00000223
    );
  blk00000003_blk000008ac : INV
    port map (
      I => blk00000003_sig00000088,
      O => blk00000003_sig00000205
    );
  blk00000003_blk000008ab : INV
    port map (
      I => blk00000003_sig0000008b,
      O => blk00000003_sig000001e7
    );
  blk00000003_blk000008aa : INV
    port map (
      I => blk00000003_sig0000008d,
      O => blk00000003_sig000001c9
    );
  blk00000003_blk000008a9 : LUT1
    generic map(
      INIT => X"1"
    )
    port map (
      I0 => blk00000003_sig0000008d,
      O => blk00000003_sig00000910
    );
  blk00000003_blk000008a8 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000567,
      I1 => blk00000003_sig0000015c,
      I2 => blk00000003_sig00000568,
      O => blk00000003_sig000008f4
    );
  blk00000003_blk000008a7 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000566,
      I1 => blk00000003_sig0000015b,
      I2 => blk00000003_sig00000568,
      O => blk00000003_sig000008f7
    );
  blk00000003_blk000008a6 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000565,
      I1 => blk00000003_sig0000015a,
      I2 => blk00000003_sig00000568,
      O => blk00000003_sig000008fa
    );
  blk00000003_blk000008a5 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000564,
      I1 => blk00000003_sig00000159,
      I2 => blk00000003_sig00000568,
      O => blk00000003_sig000008fd
    );
  blk00000003_blk000008a4 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000563,
      I1 => blk00000003_sig00000158,
      I2 => blk00000003_sig00000568,
      O => blk00000003_sig00000900
    );
  blk00000003_blk000008a3 : LUT3
    generic map(
      INIT => X"6A"
    )
    port map (
      I0 => blk00000003_sig00000562,
      I1 => blk00000003_sig00000157,
      I2 => blk00000003_sig00000568,
      O => blk00000003_sig0000090b
    );
  blk00000003_blk000008a2 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000549,
      I1 => blk00000003_sig0000054a,
      O => blk00000003_sig0000054d
    );
  blk00000003_blk000008a1 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000548,
      I1 => blk00000003_sig00000156,
      I2 => blk00000003_sig0000054a,
      O => blk00000003_sig00000550
    );
  blk00000003_blk000008a0 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000547,
      I1 => blk00000003_sig00000155,
      I2 => blk00000003_sig0000054a,
      O => blk00000003_sig00000553
    );
  blk00000003_blk0000089f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000546,
      I1 => blk00000003_sig00000154,
      I2 => blk00000003_sig0000054a,
      O => blk00000003_sig00000556
    );
  blk00000003_blk0000089e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000545,
      I1 => blk00000003_sig00000153,
      I2 => blk00000003_sig0000054a,
      O => blk00000003_sig00000559
    );
  blk00000003_blk0000089d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000544,
      I1 => blk00000003_sig00000152,
      I2 => blk00000003_sig0000054a,
      O => blk00000003_sig0000055c
    );
  blk00000003_blk0000089c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000096,
      I1 => blk00000003_sig00000151,
      I2 => blk00000003_sig0000054a,
      O => blk00000003_sig00000560
    );
  blk00000003_blk0000089b : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000052b,
      I1 => blk00000003_sig0000052c,
      O => blk00000003_sig0000052f
    );
  blk00000003_blk0000089a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000052a,
      I1 => blk00000003_sig00000150,
      I2 => blk00000003_sig0000052c,
      O => blk00000003_sig00000532
    );
  blk00000003_blk00000899 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000529,
      I1 => blk00000003_sig0000014f,
      I2 => blk00000003_sig0000052c,
      O => blk00000003_sig00000535
    );
  blk00000003_blk00000898 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000528,
      I1 => blk00000003_sig0000014e,
      I2 => blk00000003_sig0000052c,
      O => blk00000003_sig00000538
    );
  blk00000003_blk00000897 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000527,
      I1 => blk00000003_sig0000014d,
      I2 => blk00000003_sig0000052c,
      O => blk00000003_sig0000053b
    );
  blk00000003_blk00000896 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000526,
      I1 => blk00000003_sig0000014c,
      I2 => blk00000003_sig0000052c,
      O => blk00000003_sig0000053e
    );
  blk00000003_blk00000895 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000054,
      I1 => blk00000003_sig0000014b,
      I2 => blk00000003_sig0000052c,
      O => blk00000003_sig00000542
    );
  blk00000003_blk00000894 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000050d,
      I1 => blk00000003_sig0000050e,
      O => blk00000003_sig00000511
    );
  blk00000003_blk00000893 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000050c,
      I1 => blk00000003_sig0000014a,
      I2 => blk00000003_sig0000050e,
      O => blk00000003_sig00000514
    );
  blk00000003_blk00000892 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000050b,
      I1 => blk00000003_sig00000149,
      I2 => blk00000003_sig0000050e,
      O => blk00000003_sig00000517
    );
  blk00000003_blk00000891 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000050a,
      I1 => blk00000003_sig00000148,
      I2 => blk00000003_sig0000050e,
      O => blk00000003_sig0000051a
    );
  blk00000003_blk00000890 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000509,
      I1 => blk00000003_sig00000147,
      I2 => blk00000003_sig0000050e,
      O => blk00000003_sig0000051d
    );
  blk00000003_blk0000088f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000508,
      I1 => blk00000003_sig00000146,
      I2 => blk00000003_sig0000050e,
      O => blk00000003_sig00000520
    );
  blk00000003_blk0000088e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000058,
      I1 => blk00000003_sig00000145,
      I2 => blk00000003_sig0000050e,
      O => blk00000003_sig00000524
    );
  blk00000003_blk0000088d : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000004ef,
      I1 => blk00000003_sig000004f0,
      O => blk00000003_sig000004f3
    );
  blk00000003_blk0000088c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004ee,
      I1 => blk00000003_sig00000144,
      I2 => blk00000003_sig000004f0,
      O => blk00000003_sig000004f6
    );
  blk00000003_blk0000088b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004ed,
      I1 => blk00000003_sig00000143,
      I2 => blk00000003_sig000004f0,
      O => blk00000003_sig000004f9
    );
  blk00000003_blk0000088a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004ec,
      I1 => blk00000003_sig00000142,
      I2 => blk00000003_sig000004f0,
      O => blk00000003_sig000004fc
    );
  blk00000003_blk00000889 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004eb,
      I1 => blk00000003_sig00000141,
      I2 => blk00000003_sig000004f0,
      O => blk00000003_sig000004ff
    );
  blk00000003_blk00000888 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004ea,
      I1 => blk00000003_sig00000140,
      I2 => blk00000003_sig000004f0,
      O => blk00000003_sig00000502
    );
  blk00000003_blk00000887 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000005d,
      I1 => blk00000003_sig0000013f,
      I2 => blk00000003_sig000004f0,
      O => blk00000003_sig00000506
    );
  blk00000003_blk00000886 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000004d1,
      I1 => blk00000003_sig000004d2,
      O => blk00000003_sig000004d5
    );
  blk00000003_blk00000885 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004d0,
      I1 => blk00000003_sig0000013e,
      I2 => blk00000003_sig000004d2,
      O => blk00000003_sig000004d8
    );
  blk00000003_blk00000884 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004cf,
      I1 => blk00000003_sig0000013d,
      I2 => blk00000003_sig000004d2,
      O => blk00000003_sig000004db
    );
  blk00000003_blk00000883 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004ce,
      I1 => blk00000003_sig0000013c,
      I2 => blk00000003_sig000004d2,
      O => blk00000003_sig000004de
    );
  blk00000003_blk00000882 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004cd,
      I1 => blk00000003_sig0000013b,
      I2 => blk00000003_sig000004d2,
      O => blk00000003_sig000004e1
    );
  blk00000003_blk00000881 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004cc,
      I1 => blk00000003_sig0000013a,
      I2 => blk00000003_sig000004d2,
      O => blk00000003_sig000004e4
    );
  blk00000003_blk00000880 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000063,
      I1 => blk00000003_sig00000139,
      I2 => blk00000003_sig000004d2,
      O => blk00000003_sig000004e8
    );
  blk00000003_blk0000087f : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000004b3,
      I1 => blk00000003_sig000004b4,
      O => blk00000003_sig000004b7
    );
  blk00000003_blk0000087e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004b2,
      I1 => blk00000003_sig00000138,
      I2 => blk00000003_sig000004b4,
      O => blk00000003_sig000004ba
    );
  blk00000003_blk0000087d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004b1,
      I1 => blk00000003_sig00000137,
      I2 => blk00000003_sig000004b4,
      O => blk00000003_sig000004bd
    );
  blk00000003_blk0000087c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004b0,
      I1 => blk00000003_sig00000136,
      I2 => blk00000003_sig000004b4,
      O => blk00000003_sig000004c0
    );
  blk00000003_blk0000087b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004af,
      I1 => blk00000003_sig00000135,
      I2 => blk00000003_sig000004b4,
      O => blk00000003_sig000004c3
    );
  blk00000003_blk0000087a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000004ae,
      I1 => blk00000003_sig00000134,
      I2 => blk00000003_sig000004b4,
      O => blk00000003_sig000004c6
    );
  blk00000003_blk00000879 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000006a,
      I1 => blk00000003_sig00000133,
      I2 => blk00000003_sig000004b4,
      O => blk00000003_sig000004ca
    );
  blk00000003_blk00000878 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000495,
      I1 => blk00000003_sig00000496,
      O => blk00000003_sig00000499
    );
  blk00000003_blk00000877 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000494,
      I1 => blk00000003_sig00000132,
      I2 => blk00000003_sig00000496,
      O => blk00000003_sig0000049c
    );
  blk00000003_blk00000876 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000493,
      I1 => blk00000003_sig00000131,
      I2 => blk00000003_sig00000496,
      O => blk00000003_sig0000049f
    );
  blk00000003_blk00000875 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000492,
      I1 => blk00000003_sig00000130,
      I2 => blk00000003_sig00000496,
      O => blk00000003_sig000004a2
    );
  blk00000003_blk00000874 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000491,
      I1 => blk00000003_sig0000012f,
      I2 => blk00000003_sig00000496,
      O => blk00000003_sig000004a5
    );
  blk00000003_blk00000873 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000490,
      I1 => blk00000003_sig0000012e,
      I2 => blk00000003_sig00000496,
      O => blk00000003_sig000004a8
    );
  blk00000003_blk00000872 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000072,
      I1 => blk00000003_sig0000012d,
      I2 => blk00000003_sig00000496,
      O => blk00000003_sig000004ac
    );
  blk00000003_blk00000871 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000476,
      I1 => blk00000003_sig00000477,
      O => blk00000003_sig0000047a
    );
  blk00000003_blk00000870 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000475,
      I1 => blk00000003_sig0000012c,
      I2 => blk00000003_sig00000477,
      O => blk00000003_sig0000047d
    );
  blk00000003_blk0000086f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000474,
      I1 => blk00000003_sig0000012b,
      I2 => blk00000003_sig00000477,
      O => blk00000003_sig00000480
    );
  blk00000003_blk0000086e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000473,
      I1 => blk00000003_sig0000012a,
      I2 => blk00000003_sig00000477,
      O => blk00000003_sig00000483
    );
  blk00000003_blk0000086d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000472,
      I1 => blk00000003_sig00000129,
      I2 => blk00000003_sig00000477,
      O => blk00000003_sig00000486
    );
  blk00000003_blk0000086c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000471,
      I1 => blk00000003_sig00000128,
      I2 => blk00000003_sig00000477,
      O => blk00000003_sig00000489
    );
  blk00000003_blk0000086b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000048f,
      I1 => blk00000003_sig00000127,
      I2 => blk00000003_sig00000477,
      O => blk00000003_sig0000048d
    );
  blk00000003_blk0000086a : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000457,
      I1 => blk00000003_sig00000458,
      O => blk00000003_sig0000045b
    );
  blk00000003_blk00000869 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000456,
      I1 => blk00000003_sig00000126,
      I2 => blk00000003_sig00000458,
      O => blk00000003_sig0000045e
    );
  blk00000003_blk00000868 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000455,
      I1 => blk00000003_sig00000125,
      I2 => blk00000003_sig00000458,
      O => blk00000003_sig00000461
    );
  blk00000003_blk00000867 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000454,
      I1 => blk00000003_sig00000124,
      I2 => blk00000003_sig00000458,
      O => blk00000003_sig00000464
    );
  blk00000003_blk00000866 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000453,
      I1 => blk00000003_sig00000123,
      I2 => blk00000003_sig00000458,
      O => blk00000003_sig00000467
    );
  blk00000003_blk00000865 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000452,
      I1 => blk00000003_sig00000122,
      I2 => blk00000003_sig00000458,
      O => blk00000003_sig0000046a
    );
  blk00000003_blk00000864 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000470,
      I1 => blk00000003_sig00000121,
      I2 => blk00000003_sig00000458,
      O => blk00000003_sig0000046e
    );
  blk00000003_blk00000863 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000438,
      I1 => blk00000003_sig00000439,
      O => blk00000003_sig0000043c
    );
  blk00000003_blk00000862 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000437,
      I1 => blk00000003_sig00000120,
      I2 => blk00000003_sig00000439,
      O => blk00000003_sig0000043f
    );
  blk00000003_blk00000861 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000436,
      I1 => blk00000003_sig0000011f,
      I2 => blk00000003_sig00000439,
      O => blk00000003_sig00000442
    );
  blk00000003_blk00000860 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000435,
      I1 => blk00000003_sig0000011e,
      I2 => blk00000003_sig00000439,
      O => blk00000003_sig00000445
    );
  blk00000003_blk0000085f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000434,
      I1 => blk00000003_sig0000011d,
      I2 => blk00000003_sig00000439,
      O => blk00000003_sig00000448
    );
  blk00000003_blk0000085e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000433,
      I1 => blk00000003_sig0000011c,
      I2 => blk00000003_sig00000439,
      O => blk00000003_sig0000044b
    );
  blk00000003_blk0000085d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000451,
      I1 => blk00000003_sig0000011b,
      I2 => blk00000003_sig00000439,
      O => blk00000003_sig0000044f
    );
  blk00000003_blk0000085c : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000419,
      I1 => blk00000003_sig0000041a,
      O => blk00000003_sig0000041d
    );
  blk00000003_blk0000085b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000418,
      I1 => blk00000003_sig0000011a,
      I2 => blk00000003_sig0000041a,
      O => blk00000003_sig00000420
    );
  blk00000003_blk0000085a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000417,
      I1 => blk00000003_sig00000119,
      I2 => blk00000003_sig0000041a,
      O => blk00000003_sig00000423
    );
  blk00000003_blk00000859 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000416,
      I1 => blk00000003_sig00000118,
      I2 => blk00000003_sig0000041a,
      O => blk00000003_sig00000426
    );
  blk00000003_blk00000858 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000415,
      I1 => blk00000003_sig00000117,
      I2 => blk00000003_sig0000041a,
      O => blk00000003_sig00000429
    );
  blk00000003_blk00000857 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000414,
      I1 => blk00000003_sig00000116,
      I2 => blk00000003_sig0000041a,
      O => blk00000003_sig0000042c
    );
  blk00000003_blk00000856 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000432,
      I1 => blk00000003_sig00000115,
      I2 => blk00000003_sig0000041a,
      O => blk00000003_sig00000430
    );
  blk00000003_blk00000855 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000003fa,
      I1 => blk00000003_sig000003fb,
      O => blk00000003_sig000003fe
    );
  blk00000003_blk00000854 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003f9,
      I1 => blk00000003_sig00000114,
      I2 => blk00000003_sig000003fb,
      O => blk00000003_sig00000401
    );
  blk00000003_blk00000853 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003f8,
      I1 => blk00000003_sig00000113,
      I2 => blk00000003_sig000003fb,
      O => blk00000003_sig00000404
    );
  blk00000003_blk00000852 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003f7,
      I1 => blk00000003_sig00000112,
      I2 => blk00000003_sig000003fb,
      O => blk00000003_sig00000407
    );
  blk00000003_blk00000851 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003f6,
      I1 => blk00000003_sig00000111,
      I2 => blk00000003_sig000003fb,
      O => blk00000003_sig0000040a
    );
  blk00000003_blk00000850 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003f5,
      I1 => blk00000003_sig00000110,
      I2 => blk00000003_sig000003fb,
      O => blk00000003_sig0000040d
    );
  blk00000003_blk0000084f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000413,
      I1 => blk00000003_sig0000010f,
      I2 => blk00000003_sig000003fb,
      O => blk00000003_sig00000411
    );
  blk00000003_blk0000084e : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000003db,
      I1 => blk00000003_sig000003dc,
      O => blk00000003_sig000003df
    );
  blk00000003_blk0000084d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003da,
      I1 => blk00000003_sig0000010e,
      I2 => blk00000003_sig000003dc,
      O => blk00000003_sig000003e2
    );
  blk00000003_blk0000084c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003d9,
      I1 => blk00000003_sig0000010d,
      I2 => blk00000003_sig000003dc,
      O => blk00000003_sig000003e5
    );
  blk00000003_blk0000084b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003d8,
      I1 => blk00000003_sig0000010c,
      I2 => blk00000003_sig000003dc,
      O => blk00000003_sig000003e8
    );
  blk00000003_blk0000084a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003d7,
      I1 => blk00000003_sig0000010b,
      I2 => blk00000003_sig000003dc,
      O => blk00000003_sig000003eb
    );
  blk00000003_blk00000849 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003d6,
      I1 => blk00000003_sig0000010a,
      I2 => blk00000003_sig000003dc,
      O => blk00000003_sig000003ee
    );
  blk00000003_blk00000848 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003f4,
      I1 => blk00000003_sig00000109,
      I2 => blk00000003_sig000003dc,
      O => blk00000003_sig000003f2
    );
  blk00000003_blk00000847 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000003bc,
      I1 => blk00000003_sig000003bd,
      O => blk00000003_sig000003c0
    );
  blk00000003_blk00000846 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003bb,
      I1 => blk00000003_sig00000108,
      I2 => blk00000003_sig000003bd,
      O => blk00000003_sig000003c3
    );
  blk00000003_blk00000845 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003ba,
      I1 => blk00000003_sig00000107,
      I2 => blk00000003_sig000003bd,
      O => blk00000003_sig000003c6
    );
  blk00000003_blk00000844 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003b9,
      I1 => blk00000003_sig00000106,
      I2 => blk00000003_sig000003bd,
      O => blk00000003_sig000003c9
    );
  blk00000003_blk00000843 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003b8,
      I1 => blk00000003_sig00000105,
      I2 => blk00000003_sig000003bd,
      O => blk00000003_sig000003cc
    );
  blk00000003_blk00000842 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003b7,
      I1 => blk00000003_sig00000104,
      I2 => blk00000003_sig000003bd,
      O => blk00000003_sig000003cf
    );
  blk00000003_blk00000841 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003d5,
      I1 => blk00000003_sig00000103,
      I2 => blk00000003_sig000003bd,
      O => blk00000003_sig000003d3
    );
  blk00000003_blk00000840 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000039d,
      I1 => blk00000003_sig0000039e,
      O => blk00000003_sig000003a1
    );
  blk00000003_blk0000083f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000039c,
      I1 => blk00000003_sig00000102,
      I2 => blk00000003_sig0000039e,
      O => blk00000003_sig000003a4
    );
  blk00000003_blk0000083e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000039b,
      I1 => blk00000003_sig00000101,
      I2 => blk00000003_sig0000039e,
      O => blk00000003_sig000003a7
    );
  blk00000003_blk0000083d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000039a,
      I1 => blk00000003_sig00000100,
      I2 => blk00000003_sig0000039e,
      O => blk00000003_sig000003aa
    );
  blk00000003_blk0000083c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000399,
      I1 => blk00000003_sig000000ff,
      I2 => blk00000003_sig0000039e,
      O => blk00000003_sig000003ad
    );
  blk00000003_blk0000083b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000398,
      I1 => blk00000003_sig000000fe,
      I2 => blk00000003_sig0000039e,
      O => blk00000003_sig000003b0
    );
  blk00000003_blk0000083a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000003b6,
      I1 => blk00000003_sig000000fd,
      I2 => blk00000003_sig0000039e,
      O => blk00000003_sig000003b4
    );
  blk00000003_blk00000839 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000037e,
      I1 => blk00000003_sig0000037f,
      O => blk00000003_sig00000382
    );
  blk00000003_blk00000838 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000037d,
      I1 => blk00000003_sig000000fc,
      I2 => blk00000003_sig0000037f,
      O => blk00000003_sig00000385
    );
  blk00000003_blk00000837 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000037c,
      I1 => blk00000003_sig000000fb,
      I2 => blk00000003_sig0000037f,
      O => blk00000003_sig00000388
    );
  blk00000003_blk00000836 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000037b,
      I1 => blk00000003_sig000000fa,
      I2 => blk00000003_sig0000037f,
      O => blk00000003_sig0000038b
    );
  blk00000003_blk00000835 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000037a,
      I1 => blk00000003_sig000000f9,
      I2 => blk00000003_sig0000037f,
      O => blk00000003_sig0000038e
    );
  blk00000003_blk00000834 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000379,
      I1 => blk00000003_sig000000f8,
      I2 => blk00000003_sig0000037f,
      O => blk00000003_sig00000391
    );
  blk00000003_blk00000833 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000397,
      I1 => blk00000003_sig000000f7,
      I2 => blk00000003_sig0000037f,
      O => blk00000003_sig00000395
    );
  blk00000003_blk00000832 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000035f,
      I1 => blk00000003_sig00000360,
      O => blk00000003_sig00000363
    );
  blk00000003_blk00000831 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000035e,
      I1 => blk00000003_sig000000f6,
      I2 => blk00000003_sig00000360,
      O => blk00000003_sig00000366
    );
  blk00000003_blk00000830 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000035d,
      I1 => blk00000003_sig000000f5,
      I2 => blk00000003_sig00000360,
      O => blk00000003_sig00000369
    );
  blk00000003_blk0000082f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000035c,
      I1 => blk00000003_sig000000f4,
      I2 => blk00000003_sig00000360,
      O => blk00000003_sig0000036c
    );
  blk00000003_blk0000082e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000035b,
      I1 => blk00000003_sig000000f3,
      I2 => blk00000003_sig00000360,
      O => blk00000003_sig0000036f
    );
  blk00000003_blk0000082d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000035a,
      I1 => blk00000003_sig000000f2,
      I2 => blk00000003_sig00000360,
      O => blk00000003_sig00000372
    );
  blk00000003_blk0000082c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000378,
      I1 => blk00000003_sig000000f1,
      I2 => blk00000003_sig00000360,
      O => blk00000003_sig00000376
    );
  blk00000003_blk0000082b : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000340,
      I1 => blk00000003_sig00000341,
      O => blk00000003_sig00000344
    );
  blk00000003_blk0000082a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000033f,
      I1 => blk00000003_sig000000f0,
      I2 => blk00000003_sig00000341,
      O => blk00000003_sig00000347
    );
  blk00000003_blk00000829 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000033e,
      I1 => blk00000003_sig000000ef,
      I2 => blk00000003_sig00000341,
      O => blk00000003_sig0000034a
    );
  blk00000003_blk00000828 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000033d,
      I1 => blk00000003_sig000000ee,
      I2 => blk00000003_sig00000341,
      O => blk00000003_sig0000034d
    );
  blk00000003_blk00000827 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000033c,
      I1 => blk00000003_sig000000ed,
      I2 => blk00000003_sig00000341,
      O => blk00000003_sig00000350
    );
  blk00000003_blk00000826 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000033b,
      I1 => blk00000003_sig000000ec,
      I2 => blk00000003_sig00000341,
      O => blk00000003_sig00000353
    );
  blk00000003_blk00000825 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000359,
      I1 => blk00000003_sig000000eb,
      I2 => blk00000003_sig00000341,
      O => blk00000003_sig00000357
    );
  blk00000003_blk00000824 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000321,
      I1 => blk00000003_sig00000322,
      O => blk00000003_sig00000325
    );
  blk00000003_blk00000823 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000320,
      I1 => blk00000003_sig000000ea,
      I2 => blk00000003_sig00000322,
      O => blk00000003_sig00000328
    );
  blk00000003_blk00000822 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000031f,
      I1 => blk00000003_sig000000e9,
      I2 => blk00000003_sig00000322,
      O => blk00000003_sig0000032b
    );
  blk00000003_blk00000821 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000031e,
      I1 => blk00000003_sig000000e8,
      I2 => blk00000003_sig00000322,
      O => blk00000003_sig0000032e
    );
  blk00000003_blk00000820 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000031d,
      I1 => blk00000003_sig000000e7,
      I2 => blk00000003_sig00000322,
      O => blk00000003_sig00000331
    );
  blk00000003_blk0000081f : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000031c,
      I1 => blk00000003_sig000000e6,
      I2 => blk00000003_sig00000322,
      O => blk00000003_sig00000334
    );
  blk00000003_blk0000081e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000033a,
      I1 => blk00000003_sig000000e5,
      I2 => blk00000003_sig00000322,
      O => blk00000003_sig00000338
    );
  blk00000003_blk0000081d : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000302,
      I1 => blk00000003_sig00000303,
      O => blk00000003_sig00000306
    );
  blk00000003_blk0000081c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000301,
      I1 => blk00000003_sig000000e4,
      I2 => blk00000003_sig00000303,
      O => blk00000003_sig00000309
    );
  blk00000003_blk0000081b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000300,
      I1 => blk00000003_sig000000e3,
      I2 => blk00000003_sig00000303,
      O => blk00000003_sig0000030c
    );
  blk00000003_blk0000081a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002ff,
      I1 => blk00000003_sig000000e2,
      I2 => blk00000003_sig00000303,
      O => blk00000003_sig0000030f
    );
  blk00000003_blk00000819 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002fe,
      I1 => blk00000003_sig000000e1,
      I2 => blk00000003_sig00000303,
      O => blk00000003_sig00000312
    );
  blk00000003_blk00000818 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002fd,
      I1 => blk00000003_sig000000e0,
      I2 => blk00000003_sig00000303,
      O => blk00000003_sig00000315
    );
  blk00000003_blk00000817 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000031b,
      I1 => blk00000003_sig000000df,
      I2 => blk00000003_sig00000303,
      O => blk00000003_sig00000319
    );
  blk00000003_blk00000816 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000002e3,
      I1 => blk00000003_sig000002e4,
      O => blk00000003_sig000002e7
    );
  blk00000003_blk00000815 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002e2,
      I1 => blk00000003_sig000000de,
      I2 => blk00000003_sig000002e4,
      O => blk00000003_sig000002ea
    );
  blk00000003_blk00000814 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002e1,
      I1 => blk00000003_sig000000dd,
      I2 => blk00000003_sig000002e4,
      O => blk00000003_sig000002ed
    );
  blk00000003_blk00000813 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002e0,
      I1 => blk00000003_sig000000dc,
      I2 => blk00000003_sig000002e4,
      O => blk00000003_sig000002f0
    );
  blk00000003_blk00000812 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002df,
      I1 => blk00000003_sig000000db,
      I2 => blk00000003_sig000002e4,
      O => blk00000003_sig000002f3
    );
  blk00000003_blk00000811 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002de,
      I1 => blk00000003_sig000000da,
      I2 => blk00000003_sig000002e4,
      O => blk00000003_sig000002f6
    );
  blk00000003_blk00000810 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002fc,
      I1 => blk00000003_sig000000d9,
      I2 => blk00000003_sig000002e4,
      O => blk00000003_sig000002fa
    );
  blk00000003_blk0000080f : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000002c4,
      I1 => blk00000003_sig000002c5,
      O => blk00000003_sig000002c8
    );
  blk00000003_blk0000080e : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002c3,
      I1 => blk00000003_sig000000d8,
      I2 => blk00000003_sig000002c5,
      O => blk00000003_sig000002cb
    );
  blk00000003_blk0000080d : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002c2,
      I1 => blk00000003_sig000000d7,
      I2 => blk00000003_sig000002c5,
      O => blk00000003_sig000002ce
    );
  blk00000003_blk0000080c : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002c1,
      I1 => blk00000003_sig000000d6,
      I2 => blk00000003_sig000002c5,
      O => blk00000003_sig000002d1
    );
  blk00000003_blk0000080b : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002c0,
      I1 => blk00000003_sig000000d5,
      I2 => blk00000003_sig000002c5,
      O => blk00000003_sig000002d4
    );
  blk00000003_blk0000080a : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002bf,
      I1 => blk00000003_sig000000d4,
      I2 => blk00000003_sig000002c5,
      O => blk00000003_sig000002d7
    );
  blk00000003_blk00000809 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002dd,
      I1 => blk00000003_sig000000d3,
      I2 => blk00000003_sig000002c5,
      O => blk00000003_sig000002db
    );
  blk00000003_blk00000808 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000002a5,
      I1 => blk00000003_sig000002a6,
      O => blk00000003_sig000002a9
    );
  blk00000003_blk00000807 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002a4,
      I1 => blk00000003_sig000000d2,
      I2 => blk00000003_sig000002a6,
      O => blk00000003_sig000002ac
    );
  blk00000003_blk00000806 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002a3,
      I1 => blk00000003_sig000000d1,
      I2 => blk00000003_sig000002a6,
      O => blk00000003_sig000002af
    );
  blk00000003_blk00000805 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002a2,
      I1 => blk00000003_sig000000d0,
      I2 => blk00000003_sig000002a6,
      O => blk00000003_sig000002b2
    );
  blk00000003_blk00000804 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002a1,
      I1 => blk00000003_sig000000cf,
      I2 => blk00000003_sig000002a6,
      O => blk00000003_sig000002b5
    );
  blk00000003_blk00000803 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002a0,
      I1 => blk00000003_sig000000ce,
      I2 => blk00000003_sig000002a6,
      O => blk00000003_sig000002b8
    );
  blk00000003_blk00000802 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000002be,
      I1 => blk00000003_sig000000cd,
      I2 => blk00000003_sig000002a6,
      O => blk00000003_sig000002bc
    );
  blk00000003_blk00000801 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000286,
      I1 => blk00000003_sig00000287,
      O => blk00000003_sig0000028a
    );
  blk00000003_blk00000800 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000285,
      I1 => blk00000003_sig000000cc,
      I2 => blk00000003_sig00000287,
      O => blk00000003_sig0000028d
    );
  blk00000003_blk000007ff : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000284,
      I1 => blk00000003_sig000000cb,
      I2 => blk00000003_sig00000287,
      O => blk00000003_sig00000290
    );
  blk00000003_blk000007fe : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000283,
      I1 => blk00000003_sig000000ca,
      I2 => blk00000003_sig00000287,
      O => blk00000003_sig00000293
    );
  blk00000003_blk000007fd : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000282,
      I1 => blk00000003_sig000000c9,
      I2 => blk00000003_sig00000287,
      O => blk00000003_sig00000296
    );
  blk00000003_blk000007fc : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000281,
      I1 => blk00000003_sig000000c8,
      I2 => blk00000003_sig00000287,
      O => blk00000003_sig00000299
    );
  blk00000003_blk000007fb : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000029f,
      I1 => blk00000003_sig000000c7,
      I2 => blk00000003_sig00000287,
      O => blk00000003_sig0000029d
    );
  blk00000003_blk000007fa : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig00000268,
      I1 => blk00000003_sig0000008e,
      O => blk00000003_sig0000026b
    );
  blk00000003_blk000007f9 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000267,
      I1 => blk00000003_sig000000c6,
      I2 => blk00000003_sig0000008e,
      O => blk00000003_sig0000026e
    );
  blk00000003_blk000007f8 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000266,
      I1 => blk00000003_sig000000c5,
      I2 => blk00000003_sig0000008e,
      O => blk00000003_sig00000271
    );
  blk00000003_blk000007f7 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000265,
      I1 => blk00000003_sig000000c4,
      I2 => blk00000003_sig0000008e,
      O => blk00000003_sig00000274
    );
  blk00000003_blk000007f6 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000264,
      I1 => blk00000003_sig000000c3,
      I2 => blk00000003_sig0000008e,
      O => blk00000003_sig00000277
    );
  blk00000003_blk000007f5 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000263,
      I1 => blk00000003_sig000000c2,
      I2 => blk00000003_sig0000008e,
      O => blk00000003_sig0000027a
    );
  blk00000003_blk000007f4 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000280,
      I1 => blk00000003_sig000000c1,
      I2 => blk00000003_sig0000008e,
      O => blk00000003_sig0000027e
    );
  blk00000003_blk000007f3 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000024a,
      I1 => blk00000003_sig00000073,
      O => blk00000003_sig0000024d
    );
  blk00000003_blk000007f2 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000249,
      I1 => blk00000003_sig000000c0,
      I2 => blk00000003_sig00000073,
      O => blk00000003_sig00000250
    );
  blk00000003_blk000007f1 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000248,
      I1 => blk00000003_sig000000bf,
      I2 => blk00000003_sig00000073,
      O => blk00000003_sig00000253
    );
  blk00000003_blk000007f0 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000247,
      I1 => blk00000003_sig000000be,
      I2 => blk00000003_sig00000073,
      O => blk00000003_sig00000256
    );
  blk00000003_blk000007ef : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000246,
      I1 => blk00000003_sig000000bd,
      I2 => blk00000003_sig00000073,
      O => blk00000003_sig00000259
    );
  blk00000003_blk000007ee : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000245,
      I1 => blk00000003_sig000000bc,
      I2 => blk00000003_sig00000073,
      O => blk00000003_sig0000025c
    );
  blk00000003_blk000007ed : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000262,
      I1 => blk00000003_sig000000bb,
      I2 => blk00000003_sig00000073,
      O => blk00000003_sig00000260
    );
  blk00000003_blk000007ec : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000022c,
      I1 => blk00000003_sig0000007f,
      O => blk00000003_sig0000022f
    );
  blk00000003_blk000007eb : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000022b,
      I1 => blk00000003_sig000000ba,
      I2 => blk00000003_sig0000007f,
      O => blk00000003_sig00000232
    );
  blk00000003_blk000007ea : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000022a,
      I1 => blk00000003_sig000000b9,
      I2 => blk00000003_sig0000007f,
      O => blk00000003_sig00000235
    );
  blk00000003_blk000007e9 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000229,
      I1 => blk00000003_sig000000b8,
      I2 => blk00000003_sig0000007f,
      O => blk00000003_sig00000238
    );
  blk00000003_blk000007e8 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000228,
      I1 => blk00000003_sig000000b7,
      I2 => blk00000003_sig0000007f,
      O => blk00000003_sig0000023b
    );
  blk00000003_blk000007e7 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000227,
      I1 => blk00000003_sig000000b6,
      I2 => blk00000003_sig0000007f,
      O => blk00000003_sig0000023e
    );
  blk00000003_blk000007e6 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000244,
      I1 => blk00000003_sig000000b5,
      I2 => blk00000003_sig0000007f,
      O => blk00000003_sig00000242
    );
  blk00000003_blk000007e5 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000020e,
      I1 => blk00000003_sig00000084,
      O => blk00000003_sig00000211
    );
  blk00000003_blk000007e4 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000020d,
      I1 => blk00000003_sig000000b4,
      I2 => blk00000003_sig00000084,
      O => blk00000003_sig00000214
    );
  blk00000003_blk000007e3 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000020c,
      I1 => blk00000003_sig000000b3,
      I2 => blk00000003_sig00000084,
      O => blk00000003_sig00000217
    );
  blk00000003_blk000007e2 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000020b,
      I1 => blk00000003_sig000000b2,
      I2 => blk00000003_sig00000084,
      O => blk00000003_sig0000021a
    );
  blk00000003_blk000007e1 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig0000020a,
      I1 => blk00000003_sig000000b1,
      I2 => blk00000003_sig00000084,
      O => blk00000003_sig0000021d
    );
  blk00000003_blk000007e0 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000209,
      I1 => blk00000003_sig000000b0,
      I2 => blk00000003_sig00000084,
      O => blk00000003_sig00000220
    );
  blk00000003_blk000007df : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000226,
      I1 => blk00000003_sig000000af,
      I2 => blk00000003_sig00000084,
      O => blk00000003_sig00000224
    );
  blk00000003_blk000007de : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000001f0,
      I1 => blk00000003_sig00000088,
      O => blk00000003_sig000001f3
    );
  blk00000003_blk000007dd : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001ef,
      I1 => blk00000003_sig000000ae,
      I2 => blk00000003_sig00000088,
      O => blk00000003_sig000001f6
    );
  blk00000003_blk000007dc : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001ee,
      I1 => blk00000003_sig000000ad,
      I2 => blk00000003_sig00000088,
      O => blk00000003_sig000001f9
    );
  blk00000003_blk000007db : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001ed,
      I1 => blk00000003_sig000000ac,
      I2 => blk00000003_sig00000088,
      O => blk00000003_sig000001fc
    );
  blk00000003_blk000007da : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001ec,
      I1 => blk00000003_sig000000ab,
      I2 => blk00000003_sig00000088,
      O => blk00000003_sig000001ff
    );
  blk00000003_blk000007d9 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001eb,
      I1 => blk00000003_sig000000aa,
      I2 => blk00000003_sig00000088,
      O => blk00000003_sig00000202
    );
  blk00000003_blk000007d8 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig00000208,
      I1 => blk00000003_sig000000a9,
      I2 => blk00000003_sig00000088,
      O => blk00000003_sig00000206
    );
  blk00000003_blk000007d7 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000001d2,
      I1 => blk00000003_sig0000008b,
      O => blk00000003_sig000001d5
    );
  blk00000003_blk000007d6 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001d1,
      I1 => blk00000003_sig000000a8,
      I2 => blk00000003_sig0000008b,
      O => blk00000003_sig000001d8
    );
  blk00000003_blk000007d5 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001d0,
      I1 => blk00000003_sig000000a7,
      I2 => blk00000003_sig0000008b,
      O => blk00000003_sig000001db
    );
  blk00000003_blk000007d4 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001cf,
      I1 => blk00000003_sig000000a6,
      I2 => blk00000003_sig0000008b,
      O => blk00000003_sig000001de
    );
  blk00000003_blk000007d3 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001ce,
      I1 => blk00000003_sig000000a5,
      I2 => blk00000003_sig0000008b,
      O => blk00000003_sig000001e1
    );
  blk00000003_blk000007d2 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001cd,
      I1 => blk00000003_sig000000a4,
      I2 => blk00000003_sig0000008b,
      O => blk00000003_sig000001e4
    );
  blk00000003_blk000007d1 : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001ea,
      I1 => blk00000003_sig000000a3,
      I2 => blk00000003_sig0000008b,
      O => blk00000003_sig000001e8
    );
  blk00000003_blk000007d0 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig000001b5,
      I1 => blk00000003_sig0000008d,
      O => blk00000003_sig000001b7
    );
  blk00000003_blk000007cf : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001b4,
      I1 => blk00000003_sig000000a2,
      I2 => blk00000003_sig0000008d,
      O => blk00000003_sig000001ba
    );
  blk00000003_blk000007ce : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001b3,
      I1 => blk00000003_sig000000a1,
      I2 => blk00000003_sig0000008d,
      O => blk00000003_sig000001bd
    );
  blk00000003_blk000007cd : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001b2,
      I1 => blk00000003_sig000000a0,
      I2 => blk00000003_sig0000008d,
      O => blk00000003_sig000001c0
    );
  blk00000003_blk000007cc : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001b1,
      I1 => blk00000003_sig0000009f,
      I2 => blk00000003_sig0000008d,
      O => blk00000003_sig000001c3
    );
  blk00000003_blk000007cb : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001b0,
      I1 => blk00000003_sig0000009e,
      I2 => blk00000003_sig0000008d,
      O => blk00000003_sig000001c6
    );
  blk00000003_blk000007ca : LUT3
    generic map(
      INIT => X"69"
    )
    port map (
      I0 => blk00000003_sig000001cc,
      I1 => blk00000003_sig0000009d,
      I2 => blk00000003_sig0000008d,
      O => blk00000003_sig000001ca
    );
  blk00000003_blk000007c9 : LUT2
    generic map(
      INIT => X"9"
    )
    port map (
      I0 => blk00000003_sig0000017d,
      I1 => blk00000003_sig00000097,
      O => blk00000003_sig000001ae
    );
  blk00000003_blk000007c8 : LUT1
    generic map(
      INIT => X"1"
    )
    port map (
      I0 => blk00000003_sig00000568,
      O => blk00000003_sig0000017c
    );
  blk00000003_blk000007c7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000905,
      Q => blk00000003_sig0000090f
    );
  blk00000003_blk000007c6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000903,
      Q => blk00000003_sig0000090e
    );
  blk00000003_blk000007c5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008f5,
      Q => fractional(5)
    );
  blk00000003_blk000007c4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008f8,
      Q => fractional(4)
    );
  blk00000003_blk000007c3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008fb,
      Q => fractional(3)
    );
  blk00000003_blk000007c2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008fe,
      Q => fractional(2)
    );
  blk00000003_blk000007c1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000901,
      Q => fractional(1)
    );
  blk00000003_blk000007c0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000090c,
      Q => fractional(0)
    );
  blk00000003_blk000007bf : MULT_AND
    port map (
      I0 => blk00000003_sig00000157,
      I1 => blk00000003_sig00000568,
      LO => blk00000003_sig0000090d
    );
  blk00000003_blk000007be : MULT_AND
    port map (
      I0 => blk00000003_sig00000158,
      I1 => blk00000003_sig00000568,
      LO => blk00000003_sig0000090a
    );
  blk00000003_blk000007bd : MULT_AND
    port map (
      I0 => blk00000003_sig00000159,
      I1 => blk00000003_sig00000568,
      LO => blk00000003_sig00000909
    );
  blk00000003_blk000007bc : MULT_AND
    port map (
      I0 => blk00000003_sig0000015a,
      I1 => blk00000003_sig00000568,
      LO => blk00000003_sig00000908
    );
  blk00000003_blk000007bb : MULT_AND
    port map (
      I0 => blk00000003_sig0000015b,
      I1 => blk00000003_sig00000568,
      LO => blk00000003_sig00000907
    );
  blk00000003_blk000007ba : MULT_AND
    port map (
      I0 => blk00000003_sig0000015c,
      I1 => blk00000003_sig00000568,
      LO => blk00000003_sig00000906
    );
  blk00000003_blk000007b9 : MULT_AND
    port map (
      I0 => blk00000003_sig0000004f,
      I1 => blk00000003_sig00000568,
      LO => blk00000003_sig00000904
    );
  blk00000003_blk000007b8 : MUXCY
    port map (
      CI => blk00000003_sig0000004f,
      DI => blk00000003_sig0000090d,
      S => blk00000003_sig0000090b,
      O => blk00000003_sig000008ff
    );
  blk00000003_blk000007b7 : XORCY
    port map (
      CI => blk00000003_sig0000004f,
      LI => blk00000003_sig0000090b,
      O => blk00000003_sig0000090c
    );
  blk00000003_blk000007b6 : MUXCY
    port map (
      CI => blk00000003_sig000008ff,
      DI => blk00000003_sig0000090a,
      S => blk00000003_sig00000900,
      O => blk00000003_sig000008fc
    );
  blk00000003_blk000007b5 : MUXCY
    port map (
      CI => blk00000003_sig000008fc,
      DI => blk00000003_sig00000909,
      S => blk00000003_sig000008fd,
      O => blk00000003_sig000008f9
    );
  blk00000003_blk000007b4 : MUXCY
    port map (
      CI => blk00000003_sig000008f9,
      DI => blk00000003_sig00000908,
      S => blk00000003_sig000008fa,
      O => blk00000003_sig000008f6
    );
  blk00000003_blk000007b3 : MUXCY
    port map (
      CI => blk00000003_sig000008f6,
      DI => blk00000003_sig00000907,
      S => blk00000003_sig000008f7,
      O => blk00000003_sig000008f3
    );
  blk00000003_blk000007b2 : MUXCY
    port map (
      CI => blk00000003_sig000008f3,
      DI => blk00000003_sig00000906,
      S => blk00000003_sig000008f4,
      O => blk00000003_sig00000902
    );
  blk00000003_blk000007b1 : MUXCY
    port map (
      CI => blk00000003_sig00000902,
      DI => blk00000003_sig00000904,
      S => blk00000003_sig0000004f,
      O => blk00000003_sig00000905
    );
  blk00000003_blk000007b0 : XORCY
    port map (
      CI => blk00000003_sig00000902,
      LI => blk00000003_sig0000004f,
      O => blk00000003_sig00000903
    );
  blk00000003_blk000007af : XORCY
    port map (
      CI => blk00000003_sig000008ff,
      LI => blk00000003_sig00000900,
      O => blk00000003_sig00000901
    );
  blk00000003_blk000007ae : XORCY
    port map (
      CI => blk00000003_sig000008fc,
      LI => blk00000003_sig000008fd,
      O => blk00000003_sig000008fe
    );
  blk00000003_blk000007ad : XORCY
    port map (
      CI => blk00000003_sig000008f9,
      LI => blk00000003_sig000008fa,
      O => blk00000003_sig000008fb
    );
  blk00000003_blk000007ac : XORCY
    port map (
      CI => blk00000003_sig000008f6,
      LI => blk00000003_sig000008f7,
      O => blk00000003_sig000008f8
    );
  blk00000003_blk000007ab : XORCY
    port map (
      CI => blk00000003_sig000008f3,
      LI => blk00000003_sig000008f4,
      O => blk00000003_sig000008f5
    );
  blk00000003_blk000007aa : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000054a,
      Q => blk00000003_sig000008f2
    );
  blk00000003_blk000007a9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008d3,
      Q => blk00000003_sig000008f1
    );
  blk00000003_blk000007a8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008d2,
      Q => blk00000003_sig000008f0
    );
  blk00000003_blk000007a7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008d1,
      Q => blk00000003_sig000008ef
    );
  blk00000003_blk000007a6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008d0,
      Q => blk00000003_sig000008ee
    );
  blk00000003_blk000007a5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008cf,
      Q => blk00000003_sig000008ed
    );
  blk00000003_blk000007a4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008ce,
      Q => blk00000003_sig000008ec
    );
  blk00000003_blk000007a3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008cd,
      Q => blk00000003_sig000008eb
    );
  blk00000003_blk000007a2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008cc,
      Q => blk00000003_sig000008ea
    );
  blk00000003_blk000007a1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008cb,
      Q => blk00000003_sig000008e9
    );
  blk00000003_blk000007a0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008ca,
      Q => blk00000003_sig000008e8
    );
  blk00000003_blk0000079f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008c9,
      Q => blk00000003_sig000008e7
    );
  blk00000003_blk0000079e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008c8,
      Q => blk00000003_sig000008e6
    );
  blk00000003_blk0000079d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008c7,
      Q => blk00000003_sig000008e5
    );
  blk00000003_blk0000079c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008c6,
      Q => blk00000003_sig000008e4
    );
  blk00000003_blk0000079b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008c5,
      Q => blk00000003_sig000008e3
    );
  blk00000003_blk0000079a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008c4,
      Q => blk00000003_sig000008e2
    );
  blk00000003_blk00000799 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008c3,
      Q => blk00000003_sig000008e1
    );
  blk00000003_blk00000798 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008c2,
      Q => blk00000003_sig000008e0
    );
  blk00000003_blk00000797 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008c1,
      Q => blk00000003_sig000008df
    );
  blk00000003_blk00000796 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008c0,
      Q => blk00000003_sig000008de
    );
  blk00000003_blk00000795 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008bf,
      Q => blk00000003_sig000008dd
    );
  blk00000003_blk00000794 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008be,
      Q => blk00000003_sig000008dc
    );
  blk00000003_blk00000793 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008bd,
      Q => blk00000003_sig000008db
    );
  blk00000003_blk00000792 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008bc,
      Q => blk00000003_sig000008da
    );
  blk00000003_blk00000791 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008bb,
      Q => blk00000003_sig000008d9
    );
  blk00000003_blk00000790 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008ba,
      Q => blk00000003_sig000008d8
    );
  blk00000003_blk0000078f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008b9,
      Q => blk00000003_sig000008d7
    );
  blk00000003_blk0000078e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008b8,
      Q => blk00000003_sig000008d6
    );
  blk00000003_blk0000078d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008b7,
      Q => blk00000003_sig000008d5
    );
  blk00000003_blk0000078c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008b6,
      Q => blk00000003_sig000008d4
    );
  blk00000003_blk0000078b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000052c,
      Q => blk00000003_sig000008d3
    );
  blk00000003_blk0000078a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008b5,
      Q => blk00000003_sig000008d2
    );
  blk00000003_blk00000789 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008b4,
      Q => blk00000003_sig000008d1
    );
  blk00000003_blk00000788 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008b3,
      Q => blk00000003_sig000008d0
    );
  blk00000003_blk00000787 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008b2,
      Q => blk00000003_sig000008cf
    );
  blk00000003_blk00000786 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008b1,
      Q => blk00000003_sig000008ce
    );
  blk00000003_blk00000785 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008b0,
      Q => blk00000003_sig000008cd
    );
  blk00000003_blk00000784 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008af,
      Q => blk00000003_sig000008cc
    );
  blk00000003_blk00000783 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008ae,
      Q => blk00000003_sig000008cb
    );
  blk00000003_blk00000782 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008ad,
      Q => blk00000003_sig000008ca
    );
  blk00000003_blk00000781 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008ac,
      Q => blk00000003_sig000008c9
    );
  blk00000003_blk00000780 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008ab,
      Q => blk00000003_sig000008c8
    );
  blk00000003_blk0000077f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008aa,
      Q => blk00000003_sig000008c7
    );
  blk00000003_blk0000077e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008a9,
      Q => blk00000003_sig000008c6
    );
  blk00000003_blk0000077d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008a8,
      Q => blk00000003_sig000008c5
    );
  blk00000003_blk0000077c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008a7,
      Q => blk00000003_sig000008c4
    );
  blk00000003_blk0000077b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008a6,
      Q => blk00000003_sig000008c3
    );
  blk00000003_blk0000077a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008a5,
      Q => blk00000003_sig000008c2
    );
  blk00000003_blk00000779 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008a4,
      Q => blk00000003_sig000008c1
    );
  blk00000003_blk00000778 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008a3,
      Q => blk00000003_sig000008c0
    );
  blk00000003_blk00000777 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008a2,
      Q => blk00000003_sig000008bf
    );
  blk00000003_blk00000776 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008a1,
      Q => blk00000003_sig000008be
    );
  blk00000003_blk00000775 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000008a0,
      Q => blk00000003_sig000008bd
    );
  blk00000003_blk00000774 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000089f,
      Q => blk00000003_sig000008bc
    );
  blk00000003_blk00000773 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000089e,
      Q => blk00000003_sig000008bb
    );
  blk00000003_blk00000772 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000089d,
      Q => blk00000003_sig000008ba
    );
  blk00000003_blk00000771 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000089c,
      Q => blk00000003_sig000008b9
    );
  blk00000003_blk00000770 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000089b,
      Q => blk00000003_sig000008b8
    );
  blk00000003_blk0000076f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000089a,
      Q => blk00000003_sig000008b7
    );
  blk00000003_blk0000076e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000899,
      Q => blk00000003_sig000008b6
    );
  blk00000003_blk0000076d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000050e,
      Q => blk00000003_sig000008b5
    );
  blk00000003_blk0000076c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000898,
      Q => blk00000003_sig000008b4
    );
  blk00000003_blk0000076b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000897,
      Q => blk00000003_sig000008b3
    );
  blk00000003_blk0000076a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000896,
      Q => blk00000003_sig000008b2
    );
  blk00000003_blk00000769 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000895,
      Q => blk00000003_sig000008b1
    );
  blk00000003_blk00000768 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000894,
      Q => blk00000003_sig000008b0
    );
  blk00000003_blk00000767 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000893,
      Q => blk00000003_sig000008af
    );
  blk00000003_blk00000766 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000892,
      Q => blk00000003_sig000008ae
    );
  blk00000003_blk00000765 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000891,
      Q => blk00000003_sig000008ad
    );
  blk00000003_blk00000764 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000890,
      Q => blk00000003_sig000008ac
    );
  blk00000003_blk00000763 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000088f,
      Q => blk00000003_sig000008ab
    );
  blk00000003_blk00000762 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000088e,
      Q => blk00000003_sig000008aa
    );
  blk00000003_blk00000761 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000088d,
      Q => blk00000003_sig000008a9
    );
  blk00000003_blk00000760 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000088c,
      Q => blk00000003_sig000008a8
    );
  blk00000003_blk0000075f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000088b,
      Q => blk00000003_sig000008a7
    );
  blk00000003_blk0000075e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000088a,
      Q => blk00000003_sig000008a6
    );
  blk00000003_blk0000075d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000889,
      Q => blk00000003_sig000008a5
    );
  blk00000003_blk0000075c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000888,
      Q => blk00000003_sig000008a4
    );
  blk00000003_blk0000075b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000887,
      Q => blk00000003_sig000008a3
    );
  blk00000003_blk0000075a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000886,
      Q => blk00000003_sig000008a2
    );
  blk00000003_blk00000759 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000885,
      Q => blk00000003_sig000008a1
    );
  blk00000003_blk00000758 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000884,
      Q => blk00000003_sig000008a0
    );
  blk00000003_blk00000757 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000883,
      Q => blk00000003_sig0000089f
    );
  blk00000003_blk00000756 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000882,
      Q => blk00000003_sig0000089e
    );
  blk00000003_blk00000755 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000881,
      Q => blk00000003_sig0000089d
    );
  blk00000003_blk00000754 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000880,
      Q => blk00000003_sig0000089c
    );
  blk00000003_blk00000753 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000087f,
      Q => blk00000003_sig0000089b
    );
  blk00000003_blk00000752 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000087e,
      Q => blk00000003_sig0000089a
    );
  blk00000003_blk00000751 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000087d,
      Q => blk00000003_sig00000899
    );
  blk00000003_blk00000750 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004f0,
      Q => blk00000003_sig00000898
    );
  blk00000003_blk0000074f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000087c,
      Q => blk00000003_sig00000897
    );
  blk00000003_blk0000074e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000087b,
      Q => blk00000003_sig00000896
    );
  blk00000003_blk0000074d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000087a,
      Q => blk00000003_sig00000895
    );
  blk00000003_blk0000074c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000879,
      Q => blk00000003_sig00000894
    );
  blk00000003_blk0000074b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000878,
      Q => blk00000003_sig00000893
    );
  blk00000003_blk0000074a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000877,
      Q => blk00000003_sig00000892
    );
  blk00000003_blk00000749 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000876,
      Q => blk00000003_sig00000891
    );
  blk00000003_blk00000748 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000875,
      Q => blk00000003_sig00000890
    );
  blk00000003_blk00000747 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000874,
      Q => blk00000003_sig0000088f
    );
  blk00000003_blk00000746 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000873,
      Q => blk00000003_sig0000088e
    );
  blk00000003_blk00000745 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000872,
      Q => blk00000003_sig0000088d
    );
  blk00000003_blk00000744 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000871,
      Q => blk00000003_sig0000088c
    );
  blk00000003_blk00000743 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000870,
      Q => blk00000003_sig0000088b
    );
  blk00000003_blk00000742 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000086f,
      Q => blk00000003_sig0000088a
    );
  blk00000003_blk00000741 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000086e,
      Q => blk00000003_sig00000889
    );
  blk00000003_blk00000740 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000086d,
      Q => blk00000003_sig00000888
    );
  blk00000003_blk0000073f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000086c,
      Q => blk00000003_sig00000887
    );
  blk00000003_blk0000073e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000086b,
      Q => blk00000003_sig00000886
    );
  blk00000003_blk0000073d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000086a,
      Q => blk00000003_sig00000885
    );
  blk00000003_blk0000073c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000869,
      Q => blk00000003_sig00000884
    );
  blk00000003_blk0000073b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000868,
      Q => blk00000003_sig00000883
    );
  blk00000003_blk0000073a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000867,
      Q => blk00000003_sig00000882
    );
  blk00000003_blk00000739 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000866,
      Q => blk00000003_sig00000881
    );
  blk00000003_blk00000738 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000865,
      Q => blk00000003_sig00000880
    );
  blk00000003_blk00000737 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000864,
      Q => blk00000003_sig0000087f
    );
  blk00000003_blk00000736 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000863,
      Q => blk00000003_sig0000087e
    );
  blk00000003_blk00000735 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000862,
      Q => blk00000003_sig0000087d
    );
  blk00000003_blk00000734 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004d2,
      Q => blk00000003_sig0000087c
    );
  blk00000003_blk00000733 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000861,
      Q => blk00000003_sig0000087b
    );
  blk00000003_blk00000732 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000860,
      Q => blk00000003_sig0000087a
    );
  blk00000003_blk00000731 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000085f,
      Q => blk00000003_sig00000879
    );
  blk00000003_blk00000730 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000085e,
      Q => blk00000003_sig00000878
    );
  blk00000003_blk0000072f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000085d,
      Q => blk00000003_sig00000877
    );
  blk00000003_blk0000072e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000085c,
      Q => blk00000003_sig00000876
    );
  blk00000003_blk0000072d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000085b,
      Q => blk00000003_sig00000875
    );
  blk00000003_blk0000072c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000085a,
      Q => blk00000003_sig00000874
    );
  blk00000003_blk0000072b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000859,
      Q => blk00000003_sig00000873
    );
  blk00000003_blk0000072a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000858,
      Q => blk00000003_sig00000872
    );
  blk00000003_blk00000729 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000857,
      Q => blk00000003_sig00000871
    );
  blk00000003_blk00000728 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000856,
      Q => blk00000003_sig00000870
    );
  blk00000003_blk00000727 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000855,
      Q => blk00000003_sig0000086f
    );
  blk00000003_blk00000726 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000854,
      Q => blk00000003_sig0000086e
    );
  blk00000003_blk00000725 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000853,
      Q => blk00000003_sig0000086d
    );
  blk00000003_blk00000724 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000852,
      Q => blk00000003_sig0000086c
    );
  blk00000003_blk00000723 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000851,
      Q => blk00000003_sig0000086b
    );
  blk00000003_blk00000722 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000850,
      Q => blk00000003_sig0000086a
    );
  blk00000003_blk00000721 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000084f,
      Q => blk00000003_sig00000869
    );
  blk00000003_blk00000720 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000084e,
      Q => blk00000003_sig00000868
    );
  blk00000003_blk0000071f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000084d,
      Q => blk00000003_sig00000867
    );
  blk00000003_blk0000071e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000084c,
      Q => blk00000003_sig00000866
    );
  blk00000003_blk0000071d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000084b,
      Q => blk00000003_sig00000865
    );
  blk00000003_blk0000071c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000084a,
      Q => blk00000003_sig00000864
    );
  blk00000003_blk0000071b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000849,
      Q => blk00000003_sig00000863
    );
  blk00000003_blk0000071a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000848,
      Q => blk00000003_sig00000862
    );
  blk00000003_blk00000719 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004b4,
      Q => blk00000003_sig00000861
    );
  blk00000003_blk00000718 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000847,
      Q => blk00000003_sig00000860
    );
  blk00000003_blk00000717 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000846,
      Q => blk00000003_sig0000085f
    );
  blk00000003_blk00000716 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000845,
      Q => blk00000003_sig0000085e
    );
  blk00000003_blk00000715 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000844,
      Q => blk00000003_sig0000085d
    );
  blk00000003_blk00000714 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000843,
      Q => blk00000003_sig0000085c
    );
  blk00000003_blk00000713 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000842,
      Q => blk00000003_sig0000085b
    );
  blk00000003_blk00000712 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000841,
      Q => blk00000003_sig0000085a
    );
  blk00000003_blk00000711 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000840,
      Q => blk00000003_sig00000859
    );
  blk00000003_blk00000710 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000083f,
      Q => blk00000003_sig00000858
    );
  blk00000003_blk0000070f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000083e,
      Q => blk00000003_sig00000857
    );
  blk00000003_blk0000070e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000083d,
      Q => blk00000003_sig00000856
    );
  blk00000003_blk0000070d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000083c,
      Q => blk00000003_sig00000855
    );
  blk00000003_blk0000070c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000083b,
      Q => blk00000003_sig00000854
    );
  blk00000003_blk0000070b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000083a,
      Q => blk00000003_sig00000853
    );
  blk00000003_blk0000070a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000839,
      Q => blk00000003_sig00000852
    );
  blk00000003_blk00000709 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000838,
      Q => blk00000003_sig00000851
    );
  blk00000003_blk00000708 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000837,
      Q => blk00000003_sig00000850
    );
  blk00000003_blk00000707 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000836,
      Q => blk00000003_sig0000084f
    );
  blk00000003_blk00000706 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000835,
      Q => blk00000003_sig0000084e
    );
  blk00000003_blk00000705 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000834,
      Q => blk00000003_sig0000084d
    );
  blk00000003_blk00000704 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000833,
      Q => blk00000003_sig0000084c
    );
  blk00000003_blk00000703 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000832,
      Q => blk00000003_sig0000084b
    );
  blk00000003_blk00000702 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000831,
      Q => blk00000003_sig0000084a
    );
  blk00000003_blk00000701 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000830,
      Q => blk00000003_sig00000849
    );
  blk00000003_blk00000700 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000082f,
      Q => blk00000003_sig00000848
    );
  blk00000003_blk000006ff : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000496,
      Q => blk00000003_sig00000847
    );
  blk00000003_blk000006fe : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000082e,
      Q => blk00000003_sig00000846
    );
  blk00000003_blk000006fd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000082d,
      Q => blk00000003_sig00000845
    );
  blk00000003_blk000006fc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000082c,
      Q => blk00000003_sig00000844
    );
  blk00000003_blk000006fb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000082b,
      Q => blk00000003_sig00000843
    );
  blk00000003_blk000006fa : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000082a,
      Q => blk00000003_sig00000842
    );
  blk00000003_blk000006f9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000829,
      Q => blk00000003_sig00000841
    );
  blk00000003_blk000006f8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000828,
      Q => blk00000003_sig00000840
    );
  blk00000003_blk000006f7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000827,
      Q => blk00000003_sig0000083f
    );
  blk00000003_blk000006f6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000826,
      Q => blk00000003_sig0000083e
    );
  blk00000003_blk000006f5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000825,
      Q => blk00000003_sig0000083d
    );
  blk00000003_blk000006f4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000824,
      Q => blk00000003_sig0000083c
    );
  blk00000003_blk000006f3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000823,
      Q => blk00000003_sig0000083b
    );
  blk00000003_blk000006f2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000822,
      Q => blk00000003_sig0000083a
    );
  blk00000003_blk000006f1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000821,
      Q => blk00000003_sig00000839
    );
  blk00000003_blk000006f0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000820,
      Q => blk00000003_sig00000838
    );
  blk00000003_blk000006ef : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000081f,
      Q => blk00000003_sig00000837
    );
  blk00000003_blk000006ee : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000081e,
      Q => blk00000003_sig00000836
    );
  blk00000003_blk000006ed : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000081d,
      Q => blk00000003_sig00000835
    );
  blk00000003_blk000006ec : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000081c,
      Q => blk00000003_sig00000834
    );
  blk00000003_blk000006eb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000081b,
      Q => blk00000003_sig00000833
    );
  blk00000003_blk000006ea : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000081a,
      Q => blk00000003_sig00000832
    );
  blk00000003_blk000006e9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000819,
      Q => blk00000003_sig00000831
    );
  blk00000003_blk000006e8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000818,
      Q => blk00000003_sig00000830
    );
  blk00000003_blk000006e7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000817,
      Q => blk00000003_sig0000082f
    );
  blk00000003_blk000006e6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000477,
      Q => blk00000003_sig0000082e
    );
  blk00000003_blk000006e5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000816,
      Q => blk00000003_sig0000082d
    );
  blk00000003_blk000006e4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000815,
      Q => blk00000003_sig0000082c
    );
  blk00000003_blk000006e3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000814,
      Q => blk00000003_sig0000082b
    );
  blk00000003_blk000006e2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000813,
      Q => blk00000003_sig0000082a
    );
  blk00000003_blk000006e1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000812,
      Q => blk00000003_sig00000829
    );
  blk00000003_blk000006e0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000811,
      Q => blk00000003_sig00000828
    );
  blk00000003_blk000006df : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000810,
      Q => blk00000003_sig00000827
    );
  blk00000003_blk000006de : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000080f,
      Q => blk00000003_sig00000826
    );
  blk00000003_blk000006dd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000080e,
      Q => blk00000003_sig00000825
    );
  blk00000003_blk000006dc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000080d,
      Q => blk00000003_sig00000824
    );
  blk00000003_blk000006db : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000080c,
      Q => blk00000003_sig00000823
    );
  blk00000003_blk000006da : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000080b,
      Q => blk00000003_sig00000822
    );
  blk00000003_blk000006d9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000080a,
      Q => blk00000003_sig00000821
    );
  blk00000003_blk000006d8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000809,
      Q => blk00000003_sig00000820
    );
  blk00000003_blk000006d7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000808,
      Q => blk00000003_sig0000081f
    );
  blk00000003_blk000006d6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000807,
      Q => blk00000003_sig0000081e
    );
  blk00000003_blk000006d5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000806,
      Q => blk00000003_sig0000081d
    );
  blk00000003_blk000006d4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000805,
      Q => blk00000003_sig0000081c
    );
  blk00000003_blk000006d3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000804,
      Q => blk00000003_sig0000081b
    );
  blk00000003_blk000006d2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000803,
      Q => blk00000003_sig0000081a
    );
  blk00000003_blk000006d1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000802,
      Q => blk00000003_sig00000819
    );
  blk00000003_blk000006d0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000801,
      Q => blk00000003_sig00000818
    );
  blk00000003_blk000006cf : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000800,
      Q => blk00000003_sig00000817
    );
  blk00000003_blk000006ce : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007ff,
      Q => blk00000003_sig0000006b
    );
  blk00000003_blk000006cd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007fe,
      Q => blk00000003_sig0000006c
    );
  blk00000003_blk000006cc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007fd,
      Q => blk00000003_sig0000006d
    );
  blk00000003_blk000006cb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007fc,
      Q => blk00000003_sig0000006e
    );
  blk00000003_blk000006ca : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007fb,
      Q => blk00000003_sig0000006f
    );
  blk00000003_blk000006c9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007fa,
      Q => blk00000003_sig00000070
    );
  blk00000003_blk000006c8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007f9,
      Q => blk00000003_sig00000071
    );
  blk00000003_blk000006c7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007f8,
      Q => blk00000003_sig0000048f
    );
  blk00000003_blk000006c6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000458,
      Q => blk00000003_sig00000816
    );
  blk00000003_blk000006c5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007f7,
      Q => blk00000003_sig00000815
    );
  blk00000003_blk000006c4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007f6,
      Q => blk00000003_sig00000814
    );
  blk00000003_blk000006c3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007f5,
      Q => blk00000003_sig00000813
    );
  blk00000003_blk000006c2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007f4,
      Q => blk00000003_sig00000812
    );
  blk00000003_blk000006c1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007f3,
      Q => blk00000003_sig00000811
    );
  blk00000003_blk000006c0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007f2,
      Q => blk00000003_sig00000810
    );
  blk00000003_blk000006bf : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007f1,
      Q => blk00000003_sig0000080f
    );
  blk00000003_blk000006be : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007f0,
      Q => blk00000003_sig0000080e
    );
  blk00000003_blk000006bd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007ef,
      Q => blk00000003_sig0000080d
    );
  blk00000003_blk000006bc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007ee,
      Q => blk00000003_sig0000080c
    );
  blk00000003_blk000006bb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007ed,
      Q => blk00000003_sig0000080b
    );
  blk00000003_blk000006ba : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007ec,
      Q => blk00000003_sig0000080a
    );
  blk00000003_blk000006b9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007eb,
      Q => blk00000003_sig00000809
    );
  blk00000003_blk000006b8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007ea,
      Q => blk00000003_sig00000808
    );
  blk00000003_blk000006b7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007e9,
      Q => blk00000003_sig00000807
    );
  blk00000003_blk000006b6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007e8,
      Q => blk00000003_sig00000806
    );
  blk00000003_blk000006b5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007e7,
      Q => blk00000003_sig00000805
    );
  blk00000003_blk000006b4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007e6,
      Q => blk00000003_sig00000804
    );
  blk00000003_blk000006b3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007e5,
      Q => blk00000003_sig00000803
    );
  blk00000003_blk000006b2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007e4,
      Q => blk00000003_sig00000802
    );
  blk00000003_blk000006b1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007e3,
      Q => blk00000003_sig00000801
    );
  blk00000003_blk000006b0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007e2,
      Q => blk00000003_sig00000800
    );
  blk00000003_blk000006af : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007e1,
      Q => blk00000003_sig000007ff
    );
  blk00000003_blk000006ae : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007e0,
      Q => blk00000003_sig000007fe
    );
  blk00000003_blk000006ad : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007df,
      Q => blk00000003_sig000007fd
    );
  blk00000003_blk000006ac : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007de,
      Q => blk00000003_sig000007fc
    );
  blk00000003_blk000006ab : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007dd,
      Q => blk00000003_sig000007fb
    );
  blk00000003_blk000006aa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007dc,
      Q => blk00000003_sig000007fa
    );
  blk00000003_blk000006a9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007db,
      Q => blk00000003_sig000007f9
    );
  blk00000003_blk000006a8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007da,
      Q => blk00000003_sig000007f8
    );
  blk00000003_blk000006a7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007d9,
      Q => blk00000003_sig00000470
    );
  blk00000003_blk000006a6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000439,
      Q => blk00000003_sig000007f7
    );
  blk00000003_blk000006a5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007d8,
      Q => blk00000003_sig000007f6
    );
  blk00000003_blk000006a4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007d7,
      Q => blk00000003_sig000007f5
    );
  blk00000003_blk000006a3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007d6,
      Q => blk00000003_sig000007f4
    );
  blk00000003_blk000006a2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007d5,
      Q => blk00000003_sig000007f3
    );
  blk00000003_blk000006a1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007d4,
      Q => blk00000003_sig000007f2
    );
  blk00000003_blk000006a0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007d3,
      Q => blk00000003_sig000007f1
    );
  blk00000003_blk0000069f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007d2,
      Q => blk00000003_sig000007f0
    );
  blk00000003_blk0000069e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007d1,
      Q => blk00000003_sig000007ef
    );
  blk00000003_blk0000069d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007d0,
      Q => blk00000003_sig000007ee
    );
  blk00000003_blk0000069c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007cf,
      Q => blk00000003_sig000007ed
    );
  blk00000003_blk0000069b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007ce,
      Q => blk00000003_sig000007ec
    );
  blk00000003_blk0000069a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007cd,
      Q => blk00000003_sig000007eb
    );
  blk00000003_blk00000699 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007cc,
      Q => blk00000003_sig000007ea
    );
  blk00000003_blk00000698 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007cb,
      Q => blk00000003_sig000007e9
    );
  blk00000003_blk00000697 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007ca,
      Q => blk00000003_sig000007e8
    );
  blk00000003_blk00000696 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007c9,
      Q => blk00000003_sig000007e7
    );
  blk00000003_blk00000695 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007c8,
      Q => blk00000003_sig000007e6
    );
  blk00000003_blk00000694 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007c7,
      Q => blk00000003_sig000007e5
    );
  blk00000003_blk00000693 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007c6,
      Q => blk00000003_sig000007e4
    );
  blk00000003_blk00000692 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007c5,
      Q => blk00000003_sig000007e3
    );
  blk00000003_blk00000691 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007c4,
      Q => blk00000003_sig000007e2
    );
  blk00000003_blk00000690 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007c3,
      Q => blk00000003_sig000007e1
    );
  blk00000003_blk0000068f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007c2,
      Q => blk00000003_sig000007e0
    );
  blk00000003_blk0000068e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007c1,
      Q => blk00000003_sig000007df
    );
  blk00000003_blk0000068d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007c0,
      Q => blk00000003_sig000007de
    );
  blk00000003_blk0000068c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007bf,
      Q => blk00000003_sig000007dd
    );
  blk00000003_blk0000068b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007be,
      Q => blk00000003_sig000007dc
    );
  blk00000003_blk0000068a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007bd,
      Q => blk00000003_sig000007db
    );
  blk00000003_blk00000689 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007bc,
      Q => blk00000003_sig000007da
    );
  blk00000003_blk00000688 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007bb,
      Q => blk00000003_sig000007d9
    );
  blk00000003_blk00000687 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007ba,
      Q => blk00000003_sig00000451
    );
  blk00000003_blk00000686 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000041a,
      Q => blk00000003_sig000007d8
    );
  blk00000003_blk00000685 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007b9,
      Q => blk00000003_sig000007d7
    );
  blk00000003_blk00000684 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007b8,
      Q => blk00000003_sig000007d6
    );
  blk00000003_blk00000683 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007b7,
      Q => blk00000003_sig000007d5
    );
  blk00000003_blk00000682 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007b6,
      Q => blk00000003_sig000007d4
    );
  blk00000003_blk00000681 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007b5,
      Q => blk00000003_sig000007d3
    );
  blk00000003_blk00000680 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007b4,
      Q => blk00000003_sig000007d2
    );
  blk00000003_blk0000067f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007b3,
      Q => blk00000003_sig000007d1
    );
  blk00000003_blk0000067e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007b2,
      Q => blk00000003_sig000007d0
    );
  blk00000003_blk0000067d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007b1,
      Q => blk00000003_sig000007cf
    );
  blk00000003_blk0000067c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007b0,
      Q => blk00000003_sig000007ce
    );
  blk00000003_blk0000067b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007af,
      Q => blk00000003_sig000007cd
    );
  blk00000003_blk0000067a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007ae,
      Q => blk00000003_sig000007cc
    );
  blk00000003_blk00000679 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007ad,
      Q => blk00000003_sig000007cb
    );
  blk00000003_blk00000678 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007ac,
      Q => blk00000003_sig000007ca
    );
  blk00000003_blk00000677 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007ab,
      Q => blk00000003_sig000007c9
    );
  blk00000003_blk00000676 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007aa,
      Q => blk00000003_sig000007c8
    );
  blk00000003_blk00000675 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007a9,
      Q => blk00000003_sig000007c7
    );
  blk00000003_blk00000674 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007a8,
      Q => blk00000003_sig000007c6
    );
  blk00000003_blk00000673 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007a7,
      Q => blk00000003_sig000007c5
    );
  blk00000003_blk00000672 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007a6,
      Q => blk00000003_sig000007c4
    );
  blk00000003_blk00000671 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007a5,
      Q => blk00000003_sig000007c3
    );
  blk00000003_blk00000670 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007a4,
      Q => blk00000003_sig000007c2
    );
  blk00000003_blk0000066f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007a3,
      Q => blk00000003_sig000007c1
    );
  blk00000003_blk0000066e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007a2,
      Q => blk00000003_sig000007c0
    );
  blk00000003_blk0000066d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007a1,
      Q => blk00000003_sig000007bf
    );
  blk00000003_blk0000066c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000007a0,
      Q => blk00000003_sig000007be
    );
  blk00000003_blk0000066b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000079f,
      Q => blk00000003_sig000007bd
    );
  blk00000003_blk0000066a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000079e,
      Q => blk00000003_sig000007bc
    );
  blk00000003_blk00000669 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000079d,
      Q => blk00000003_sig000007bb
    );
  blk00000003_blk00000668 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000079c,
      Q => blk00000003_sig000007ba
    );
  blk00000003_blk00000667 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000079b,
      Q => blk00000003_sig00000432
    );
  blk00000003_blk00000666 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003fb,
      Q => blk00000003_sig000007b9
    );
  blk00000003_blk00000665 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000079a,
      Q => blk00000003_sig000007b8
    );
  blk00000003_blk00000664 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000799,
      Q => blk00000003_sig000007b7
    );
  blk00000003_blk00000663 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000798,
      Q => blk00000003_sig000007b6
    );
  blk00000003_blk00000662 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000797,
      Q => blk00000003_sig000007b5
    );
  blk00000003_blk00000661 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000796,
      Q => blk00000003_sig000007b4
    );
  blk00000003_blk00000660 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000795,
      Q => blk00000003_sig000007b3
    );
  blk00000003_blk0000065f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000794,
      Q => blk00000003_sig000007b2
    );
  blk00000003_blk0000065e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000793,
      Q => blk00000003_sig000007b1
    );
  blk00000003_blk0000065d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000792,
      Q => blk00000003_sig000007b0
    );
  blk00000003_blk0000065c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000791,
      Q => blk00000003_sig000007af
    );
  blk00000003_blk0000065b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000790,
      Q => blk00000003_sig000007ae
    );
  blk00000003_blk0000065a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000078f,
      Q => blk00000003_sig000007ad
    );
  blk00000003_blk00000659 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000078e,
      Q => blk00000003_sig000007ac
    );
  blk00000003_blk00000658 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000078d,
      Q => blk00000003_sig000007ab
    );
  blk00000003_blk00000657 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000078c,
      Q => blk00000003_sig000007aa
    );
  blk00000003_blk00000656 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000078b,
      Q => blk00000003_sig000007a9
    );
  blk00000003_blk00000655 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000078a,
      Q => blk00000003_sig000007a8
    );
  blk00000003_blk00000654 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000789,
      Q => blk00000003_sig000007a7
    );
  blk00000003_blk00000653 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000788,
      Q => blk00000003_sig000007a6
    );
  blk00000003_blk00000652 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000787,
      Q => blk00000003_sig000007a5
    );
  blk00000003_blk00000651 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000786,
      Q => blk00000003_sig000007a4
    );
  blk00000003_blk00000650 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000785,
      Q => blk00000003_sig000007a3
    );
  blk00000003_blk0000064f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000784,
      Q => blk00000003_sig000007a2
    );
  blk00000003_blk0000064e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000783,
      Q => blk00000003_sig000007a1
    );
  blk00000003_blk0000064d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000782,
      Q => blk00000003_sig000007a0
    );
  blk00000003_blk0000064c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000781,
      Q => blk00000003_sig0000079f
    );
  blk00000003_blk0000064b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000780,
      Q => blk00000003_sig0000079e
    );
  blk00000003_blk0000064a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000077f,
      Q => blk00000003_sig0000079d
    );
  blk00000003_blk00000649 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000077e,
      Q => blk00000003_sig0000079c
    );
  blk00000003_blk00000648 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000077d,
      Q => blk00000003_sig0000079b
    );
  blk00000003_blk00000647 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000077c,
      Q => blk00000003_sig00000413
    );
  blk00000003_blk00000646 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003dc,
      Q => blk00000003_sig0000079a
    );
  blk00000003_blk00000645 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000077b,
      Q => blk00000003_sig00000799
    );
  blk00000003_blk00000644 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000077a,
      Q => blk00000003_sig00000798
    );
  blk00000003_blk00000643 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000779,
      Q => blk00000003_sig00000797
    );
  blk00000003_blk00000642 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000778,
      Q => blk00000003_sig00000796
    );
  blk00000003_blk00000641 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000777,
      Q => blk00000003_sig00000795
    );
  blk00000003_blk00000640 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000776,
      Q => blk00000003_sig00000794
    );
  blk00000003_blk0000063f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000775,
      Q => blk00000003_sig00000793
    );
  blk00000003_blk0000063e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000774,
      Q => blk00000003_sig00000792
    );
  blk00000003_blk0000063d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000773,
      Q => blk00000003_sig00000791
    );
  blk00000003_blk0000063c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000772,
      Q => blk00000003_sig00000790
    );
  blk00000003_blk0000063b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000771,
      Q => blk00000003_sig0000078f
    );
  blk00000003_blk0000063a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000770,
      Q => blk00000003_sig0000078e
    );
  blk00000003_blk00000639 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000076f,
      Q => blk00000003_sig0000078d
    );
  blk00000003_blk00000638 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000076e,
      Q => blk00000003_sig0000078c
    );
  blk00000003_blk00000637 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000076d,
      Q => blk00000003_sig0000078b
    );
  blk00000003_blk00000636 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000076c,
      Q => blk00000003_sig0000078a
    );
  blk00000003_blk00000635 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000076b,
      Q => blk00000003_sig00000789
    );
  blk00000003_blk00000634 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000076a,
      Q => blk00000003_sig00000788
    );
  blk00000003_blk00000633 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000769,
      Q => blk00000003_sig00000787
    );
  blk00000003_blk00000632 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000768,
      Q => blk00000003_sig00000786
    );
  blk00000003_blk00000631 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000767,
      Q => blk00000003_sig00000785
    );
  blk00000003_blk00000630 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000766,
      Q => blk00000003_sig00000784
    );
  blk00000003_blk0000062f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000765,
      Q => blk00000003_sig00000783
    );
  blk00000003_blk0000062e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000764,
      Q => blk00000003_sig00000782
    );
  blk00000003_blk0000062d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000763,
      Q => blk00000003_sig00000781
    );
  blk00000003_blk0000062c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000762,
      Q => blk00000003_sig00000780
    );
  blk00000003_blk0000062b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000761,
      Q => blk00000003_sig0000077f
    );
  blk00000003_blk0000062a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000760,
      Q => blk00000003_sig0000077e
    );
  blk00000003_blk00000629 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000075f,
      Q => blk00000003_sig0000077d
    );
  blk00000003_blk00000628 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000075e,
      Q => blk00000003_sig0000077c
    );
  blk00000003_blk00000627 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000075d,
      Q => blk00000003_sig000003f4
    );
  blk00000003_blk00000626 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003bd,
      Q => blk00000003_sig0000077b
    );
  blk00000003_blk00000625 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000075c,
      Q => blk00000003_sig0000077a
    );
  blk00000003_blk00000624 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000075b,
      Q => blk00000003_sig00000779
    );
  blk00000003_blk00000623 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000075a,
      Q => blk00000003_sig00000778
    );
  blk00000003_blk00000622 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000759,
      Q => blk00000003_sig00000777
    );
  blk00000003_blk00000621 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000758,
      Q => blk00000003_sig00000776
    );
  blk00000003_blk00000620 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000757,
      Q => blk00000003_sig00000775
    );
  blk00000003_blk0000061f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000756,
      Q => blk00000003_sig00000774
    );
  blk00000003_blk0000061e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000755,
      Q => blk00000003_sig00000773
    );
  blk00000003_blk0000061d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000754,
      Q => blk00000003_sig00000772
    );
  blk00000003_blk0000061c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000753,
      Q => blk00000003_sig00000771
    );
  blk00000003_blk0000061b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000752,
      Q => blk00000003_sig00000770
    );
  blk00000003_blk0000061a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000751,
      Q => blk00000003_sig0000076f
    );
  blk00000003_blk00000619 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000750,
      Q => blk00000003_sig0000076e
    );
  blk00000003_blk00000618 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000074f,
      Q => blk00000003_sig0000076d
    );
  blk00000003_blk00000617 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000074e,
      Q => blk00000003_sig0000076c
    );
  blk00000003_blk00000616 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000074d,
      Q => blk00000003_sig0000076b
    );
  blk00000003_blk00000615 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000074c,
      Q => blk00000003_sig0000076a
    );
  blk00000003_blk00000614 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000074b,
      Q => blk00000003_sig00000769
    );
  blk00000003_blk00000613 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000074a,
      Q => blk00000003_sig00000768
    );
  blk00000003_blk00000612 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000749,
      Q => blk00000003_sig00000767
    );
  blk00000003_blk00000611 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000748,
      Q => blk00000003_sig00000766
    );
  blk00000003_blk00000610 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000747,
      Q => blk00000003_sig00000765
    );
  blk00000003_blk0000060f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000746,
      Q => blk00000003_sig00000764
    );
  blk00000003_blk0000060e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000745,
      Q => blk00000003_sig00000763
    );
  blk00000003_blk0000060d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000744,
      Q => blk00000003_sig00000762
    );
  blk00000003_blk0000060c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000743,
      Q => blk00000003_sig00000761
    );
  blk00000003_blk0000060b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000742,
      Q => blk00000003_sig00000760
    );
  blk00000003_blk0000060a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000741,
      Q => blk00000003_sig0000075f
    );
  blk00000003_blk00000609 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000740,
      Q => blk00000003_sig0000075e
    );
  blk00000003_blk00000608 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000073f,
      Q => blk00000003_sig0000075d
    );
  blk00000003_blk00000607 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000073e,
      Q => blk00000003_sig000003d5
    );
  blk00000003_blk00000606 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000039e,
      Q => blk00000003_sig0000075c
    );
  blk00000003_blk00000605 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000073d,
      Q => blk00000003_sig0000075b
    );
  blk00000003_blk00000604 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000073c,
      Q => blk00000003_sig0000075a
    );
  blk00000003_blk00000603 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000073b,
      Q => blk00000003_sig00000759
    );
  blk00000003_blk00000602 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000073a,
      Q => blk00000003_sig00000758
    );
  blk00000003_blk00000601 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000739,
      Q => blk00000003_sig00000757
    );
  blk00000003_blk00000600 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000738,
      Q => blk00000003_sig00000756
    );
  blk00000003_blk000005ff : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000737,
      Q => blk00000003_sig00000755
    );
  blk00000003_blk000005fe : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000736,
      Q => blk00000003_sig00000754
    );
  blk00000003_blk000005fd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000735,
      Q => blk00000003_sig00000753
    );
  blk00000003_blk000005fc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000734,
      Q => blk00000003_sig00000752
    );
  blk00000003_blk000005fb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000733,
      Q => blk00000003_sig00000751
    );
  blk00000003_blk000005fa : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000732,
      Q => blk00000003_sig00000750
    );
  blk00000003_blk000005f9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000731,
      Q => blk00000003_sig0000074f
    );
  blk00000003_blk000005f8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000730,
      Q => blk00000003_sig0000074e
    );
  blk00000003_blk000005f7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000072f,
      Q => blk00000003_sig0000074d
    );
  blk00000003_blk000005f6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000072e,
      Q => blk00000003_sig0000074c
    );
  blk00000003_blk000005f5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000072d,
      Q => blk00000003_sig0000074b
    );
  blk00000003_blk000005f4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000072c,
      Q => blk00000003_sig0000074a
    );
  blk00000003_blk000005f3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000072b,
      Q => blk00000003_sig00000749
    );
  blk00000003_blk000005f2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000072a,
      Q => blk00000003_sig00000748
    );
  blk00000003_blk000005f1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000729,
      Q => blk00000003_sig00000747
    );
  blk00000003_blk000005f0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000728,
      Q => blk00000003_sig00000746
    );
  blk00000003_blk000005ef : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000727,
      Q => blk00000003_sig00000745
    );
  blk00000003_blk000005ee : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000726,
      Q => blk00000003_sig00000744
    );
  blk00000003_blk000005ed : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000725,
      Q => blk00000003_sig00000743
    );
  blk00000003_blk000005ec : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000724,
      Q => blk00000003_sig00000742
    );
  blk00000003_blk000005eb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000723,
      Q => blk00000003_sig00000741
    );
  blk00000003_blk000005ea : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000722,
      Q => blk00000003_sig00000740
    );
  blk00000003_blk000005e9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000721,
      Q => blk00000003_sig0000073f
    );
  blk00000003_blk000005e8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000720,
      Q => blk00000003_sig0000073e
    );
  blk00000003_blk000005e7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000071f,
      Q => blk00000003_sig000003b6
    );
  blk00000003_blk000005e6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000037f,
      Q => blk00000003_sig0000073d
    );
  blk00000003_blk000005e5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000071e,
      Q => blk00000003_sig0000073c
    );
  blk00000003_blk000005e4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000071d,
      Q => blk00000003_sig0000073b
    );
  blk00000003_blk000005e3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000071c,
      Q => blk00000003_sig0000073a
    );
  blk00000003_blk000005e2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000071b,
      Q => blk00000003_sig00000739
    );
  blk00000003_blk000005e1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000071a,
      Q => blk00000003_sig00000738
    );
  blk00000003_blk000005e0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000719,
      Q => blk00000003_sig00000737
    );
  blk00000003_blk000005df : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000718,
      Q => blk00000003_sig00000736
    );
  blk00000003_blk000005de : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000717,
      Q => blk00000003_sig00000735
    );
  blk00000003_blk000005dd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000716,
      Q => blk00000003_sig00000734
    );
  blk00000003_blk000005dc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000715,
      Q => blk00000003_sig00000733
    );
  blk00000003_blk000005db : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000714,
      Q => blk00000003_sig00000732
    );
  blk00000003_blk000005da : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000713,
      Q => blk00000003_sig00000731
    );
  blk00000003_blk000005d9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000712,
      Q => blk00000003_sig00000730
    );
  blk00000003_blk000005d8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000711,
      Q => blk00000003_sig0000072f
    );
  blk00000003_blk000005d7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000710,
      Q => blk00000003_sig0000072e
    );
  blk00000003_blk000005d6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000070f,
      Q => blk00000003_sig0000072d
    );
  blk00000003_blk000005d5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000070e,
      Q => blk00000003_sig0000072c
    );
  blk00000003_blk000005d4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000070d,
      Q => blk00000003_sig0000072b
    );
  blk00000003_blk000005d3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000070c,
      Q => blk00000003_sig0000072a
    );
  blk00000003_blk000005d2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000070b,
      Q => blk00000003_sig00000729
    );
  blk00000003_blk000005d1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000070a,
      Q => blk00000003_sig00000728
    );
  blk00000003_blk000005d0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000709,
      Q => blk00000003_sig00000727
    );
  blk00000003_blk000005cf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000708,
      Q => blk00000003_sig00000726
    );
  blk00000003_blk000005ce : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000707,
      Q => blk00000003_sig00000725
    );
  blk00000003_blk000005cd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000706,
      Q => blk00000003_sig00000724
    );
  blk00000003_blk000005cc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000705,
      Q => blk00000003_sig00000723
    );
  blk00000003_blk000005cb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000704,
      Q => blk00000003_sig00000722
    );
  blk00000003_blk000005ca : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000703,
      Q => blk00000003_sig00000721
    );
  blk00000003_blk000005c9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000702,
      Q => blk00000003_sig00000720
    );
  blk00000003_blk000005c8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000701,
      Q => blk00000003_sig0000071f
    );
  blk00000003_blk000005c7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000700,
      Q => blk00000003_sig00000397
    );
  blk00000003_blk000005c6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000360,
      Q => blk00000003_sig0000071e
    );
  blk00000003_blk000005c5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ff,
      Q => blk00000003_sig0000071d
    );
  blk00000003_blk000005c4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006fe,
      Q => blk00000003_sig0000071c
    );
  blk00000003_blk000005c3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006fd,
      Q => blk00000003_sig0000071b
    );
  blk00000003_blk000005c2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006fc,
      Q => blk00000003_sig0000071a
    );
  blk00000003_blk000005c1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006fb,
      Q => blk00000003_sig00000719
    );
  blk00000003_blk000005c0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006fa,
      Q => blk00000003_sig00000718
    );
  blk00000003_blk000005bf : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006f9,
      Q => blk00000003_sig00000717
    );
  blk00000003_blk000005be : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006f8,
      Q => blk00000003_sig00000716
    );
  blk00000003_blk000005bd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006f7,
      Q => blk00000003_sig00000715
    );
  blk00000003_blk000005bc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006f6,
      Q => blk00000003_sig00000714
    );
  blk00000003_blk000005bb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006f5,
      Q => blk00000003_sig00000713
    );
  blk00000003_blk000005ba : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006f4,
      Q => blk00000003_sig00000712
    );
  blk00000003_blk000005b9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006f3,
      Q => blk00000003_sig00000711
    );
  blk00000003_blk000005b8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006f2,
      Q => blk00000003_sig00000710
    );
  blk00000003_blk000005b7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006f1,
      Q => blk00000003_sig0000070f
    );
  blk00000003_blk000005b6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006f0,
      Q => blk00000003_sig0000070e
    );
  blk00000003_blk000005b5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ef,
      Q => blk00000003_sig0000070d
    );
  blk00000003_blk000005b4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ee,
      Q => blk00000003_sig0000070c
    );
  blk00000003_blk000005b3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ed,
      Q => blk00000003_sig0000070b
    );
  blk00000003_blk000005b2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ec,
      Q => blk00000003_sig0000070a
    );
  blk00000003_blk000005b1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006eb,
      Q => blk00000003_sig00000709
    );
  blk00000003_blk000005b0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ea,
      Q => blk00000003_sig00000708
    );
  blk00000003_blk000005af : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006e9,
      Q => blk00000003_sig00000707
    );
  blk00000003_blk000005ae : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006e8,
      Q => blk00000003_sig00000706
    );
  blk00000003_blk000005ad : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006e7,
      Q => blk00000003_sig00000705
    );
  blk00000003_blk000005ac : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006e6,
      Q => blk00000003_sig00000704
    );
  blk00000003_blk000005ab : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006e5,
      Q => blk00000003_sig00000703
    );
  blk00000003_blk000005aa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006e4,
      Q => blk00000003_sig00000702
    );
  blk00000003_blk000005a9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006e3,
      Q => blk00000003_sig00000701
    );
  blk00000003_blk000005a8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006e2,
      Q => blk00000003_sig00000700
    );
  blk00000003_blk000005a7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006e1,
      Q => blk00000003_sig00000378
    );
  blk00000003_blk000005a6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000341,
      Q => blk00000003_sig000006ff
    );
  blk00000003_blk000005a5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006e0,
      Q => blk00000003_sig000006fe
    );
  blk00000003_blk000005a4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006df,
      Q => blk00000003_sig000006fd
    );
  blk00000003_blk000005a3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006de,
      Q => blk00000003_sig000006fc
    );
  blk00000003_blk000005a2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006dd,
      Q => blk00000003_sig000006fb
    );
  blk00000003_blk000005a1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006dc,
      Q => blk00000003_sig000006fa
    );
  blk00000003_blk000005a0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006db,
      Q => blk00000003_sig000006f9
    );
  blk00000003_blk0000059f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006da,
      Q => blk00000003_sig000006f8
    );
  blk00000003_blk0000059e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006d9,
      Q => blk00000003_sig000006f7
    );
  blk00000003_blk0000059d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006d8,
      Q => blk00000003_sig000006f6
    );
  blk00000003_blk0000059c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006d7,
      Q => blk00000003_sig000006f5
    );
  blk00000003_blk0000059b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006d6,
      Q => blk00000003_sig000006f4
    );
  blk00000003_blk0000059a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006d5,
      Q => blk00000003_sig000006f3
    );
  blk00000003_blk00000599 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006d4,
      Q => blk00000003_sig000006f2
    );
  blk00000003_blk00000598 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006d3,
      Q => blk00000003_sig000006f1
    );
  blk00000003_blk00000597 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006d2,
      Q => blk00000003_sig000006f0
    );
  blk00000003_blk00000596 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006d1,
      Q => blk00000003_sig000006ef
    );
  blk00000003_blk00000595 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006d0,
      Q => blk00000003_sig000006ee
    );
  blk00000003_blk00000594 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006cf,
      Q => blk00000003_sig000006ed
    );
  blk00000003_blk00000593 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ce,
      Q => blk00000003_sig000006ec
    );
  blk00000003_blk00000592 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006cd,
      Q => blk00000003_sig000006eb
    );
  blk00000003_blk00000591 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006cc,
      Q => blk00000003_sig000006ea
    );
  blk00000003_blk00000590 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006cb,
      Q => blk00000003_sig000006e9
    );
  blk00000003_blk0000058f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ca,
      Q => blk00000003_sig000006e8
    );
  blk00000003_blk0000058e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006c9,
      Q => blk00000003_sig000006e7
    );
  blk00000003_blk0000058d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006c8,
      Q => blk00000003_sig000006e6
    );
  blk00000003_blk0000058c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006c7,
      Q => blk00000003_sig000006e5
    );
  blk00000003_blk0000058b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006c6,
      Q => blk00000003_sig000006e4
    );
  blk00000003_blk0000058a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006c5,
      Q => blk00000003_sig000006e3
    );
  blk00000003_blk00000589 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006c4,
      Q => blk00000003_sig000006e2
    );
  blk00000003_blk00000588 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006c3,
      Q => blk00000003_sig000006e1
    );
  blk00000003_blk00000587 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006c2,
      Q => blk00000003_sig00000359
    );
  blk00000003_blk00000586 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000322,
      Q => blk00000003_sig000006e0
    );
  blk00000003_blk00000585 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006c1,
      Q => blk00000003_sig000006df
    );
  blk00000003_blk00000584 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006c0,
      Q => blk00000003_sig000006de
    );
  blk00000003_blk00000583 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006bf,
      Q => blk00000003_sig000006dd
    );
  blk00000003_blk00000582 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006be,
      Q => blk00000003_sig000006dc
    );
  blk00000003_blk00000581 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006bd,
      Q => blk00000003_sig000006db
    );
  blk00000003_blk00000580 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006bc,
      Q => blk00000003_sig000006da
    );
  blk00000003_blk0000057f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006bb,
      Q => blk00000003_sig000006d9
    );
  blk00000003_blk0000057e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ba,
      Q => blk00000003_sig000006d8
    );
  blk00000003_blk0000057d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006b9,
      Q => blk00000003_sig000006d7
    );
  blk00000003_blk0000057c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006b8,
      Q => blk00000003_sig000006d6
    );
  blk00000003_blk0000057b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006b7,
      Q => blk00000003_sig000006d5
    );
  blk00000003_blk0000057a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006b6,
      Q => blk00000003_sig000006d4
    );
  blk00000003_blk00000579 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006b5,
      Q => blk00000003_sig000006d3
    );
  blk00000003_blk00000578 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006b4,
      Q => blk00000003_sig000006d2
    );
  blk00000003_blk00000577 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006b3,
      Q => blk00000003_sig000006d1
    );
  blk00000003_blk00000576 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006b2,
      Q => blk00000003_sig000006d0
    );
  blk00000003_blk00000575 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006b1,
      Q => blk00000003_sig000006cf
    );
  blk00000003_blk00000574 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006b0,
      Q => blk00000003_sig000006ce
    );
  blk00000003_blk00000573 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006af,
      Q => blk00000003_sig000006cd
    );
  blk00000003_blk00000572 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ae,
      Q => blk00000003_sig000006cc
    );
  blk00000003_blk00000571 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ad,
      Q => blk00000003_sig000006cb
    );
  blk00000003_blk00000570 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ac,
      Q => blk00000003_sig000006ca
    );
  blk00000003_blk0000056f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006ab,
      Q => blk00000003_sig000006c9
    );
  blk00000003_blk0000056e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006aa,
      Q => blk00000003_sig000006c8
    );
  blk00000003_blk0000056d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a9,
      Q => blk00000003_sig000006c7
    );
  blk00000003_blk0000056c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a8,
      Q => blk00000003_sig000006c6
    );
  blk00000003_blk0000056b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a7,
      Q => blk00000003_sig000006c5
    );
  blk00000003_blk0000056a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a6,
      Q => blk00000003_sig000006c4
    );
  blk00000003_blk00000569 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a5,
      Q => blk00000003_sig000006c3
    );
  blk00000003_blk00000568 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a4,
      Q => blk00000003_sig000006c2
    );
  blk00000003_blk00000567 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a3,
      Q => blk00000003_sig0000033a
    );
  blk00000003_blk00000566 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000303,
      Q => blk00000003_sig000006c1
    );
  blk00000003_blk00000565 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a2,
      Q => blk00000003_sig000006c0
    );
  blk00000003_blk00000564 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a1,
      Q => blk00000003_sig000006bf
    );
  blk00000003_blk00000563 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000006a0,
      Q => blk00000003_sig000006be
    );
  blk00000003_blk00000562 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000069f,
      Q => blk00000003_sig000006bd
    );
  blk00000003_blk00000561 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000069e,
      Q => blk00000003_sig000006bc
    );
  blk00000003_blk00000560 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000069d,
      Q => blk00000003_sig000006bb
    );
  blk00000003_blk0000055f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000069c,
      Q => blk00000003_sig000006ba
    );
  blk00000003_blk0000055e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000069b,
      Q => blk00000003_sig000006b9
    );
  blk00000003_blk0000055d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000069a,
      Q => blk00000003_sig000006b8
    );
  blk00000003_blk0000055c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000699,
      Q => blk00000003_sig000006b7
    );
  blk00000003_blk0000055b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000698,
      Q => blk00000003_sig000006b6
    );
  blk00000003_blk0000055a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000697,
      Q => blk00000003_sig000006b5
    );
  blk00000003_blk00000559 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000696,
      Q => blk00000003_sig000006b4
    );
  blk00000003_blk00000558 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000695,
      Q => blk00000003_sig000006b3
    );
  blk00000003_blk00000557 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000694,
      Q => blk00000003_sig000006b2
    );
  blk00000003_blk00000556 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000693,
      Q => blk00000003_sig000006b1
    );
  blk00000003_blk00000555 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000692,
      Q => blk00000003_sig000006b0
    );
  blk00000003_blk00000554 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000691,
      Q => blk00000003_sig000006af
    );
  blk00000003_blk00000553 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000690,
      Q => blk00000003_sig000006ae
    );
  blk00000003_blk00000552 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000068f,
      Q => blk00000003_sig000006ad
    );
  blk00000003_blk00000551 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000068e,
      Q => blk00000003_sig000006ac
    );
  blk00000003_blk00000550 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000068d,
      Q => blk00000003_sig000006ab
    );
  blk00000003_blk0000054f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000068c,
      Q => blk00000003_sig000006aa
    );
  blk00000003_blk0000054e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000068b,
      Q => blk00000003_sig000006a9
    );
  blk00000003_blk0000054d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000068a,
      Q => blk00000003_sig000006a8
    );
  blk00000003_blk0000054c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000689,
      Q => blk00000003_sig000006a7
    );
  blk00000003_blk0000054b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000688,
      Q => blk00000003_sig000006a6
    );
  blk00000003_blk0000054a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000687,
      Q => blk00000003_sig000006a5
    );
  blk00000003_blk00000549 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000686,
      Q => blk00000003_sig000006a4
    );
  blk00000003_blk00000548 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000685,
      Q => blk00000003_sig000006a3
    );
  blk00000003_blk00000547 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000684,
      Q => blk00000003_sig0000031b
    );
  blk00000003_blk00000546 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002e4,
      Q => blk00000003_sig000006a2
    );
  blk00000003_blk00000545 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000683,
      Q => blk00000003_sig000006a1
    );
  blk00000003_blk00000544 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000682,
      Q => blk00000003_sig000006a0
    );
  blk00000003_blk00000543 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000681,
      Q => blk00000003_sig0000069f
    );
  blk00000003_blk00000542 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000680,
      Q => blk00000003_sig0000069e
    );
  blk00000003_blk00000541 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000067f,
      Q => blk00000003_sig0000069d
    );
  blk00000003_blk00000540 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000067e,
      Q => blk00000003_sig0000069c
    );
  blk00000003_blk0000053f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000067d,
      Q => blk00000003_sig0000069b
    );
  blk00000003_blk0000053e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000067c,
      Q => blk00000003_sig0000069a
    );
  blk00000003_blk0000053d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000067b,
      Q => blk00000003_sig00000699
    );
  blk00000003_blk0000053c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000067a,
      Q => blk00000003_sig00000698
    );
  blk00000003_blk0000053b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000679,
      Q => blk00000003_sig00000697
    );
  blk00000003_blk0000053a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000678,
      Q => blk00000003_sig00000696
    );
  blk00000003_blk00000539 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000677,
      Q => blk00000003_sig00000695
    );
  blk00000003_blk00000538 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000676,
      Q => blk00000003_sig00000694
    );
  blk00000003_blk00000537 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000675,
      Q => blk00000003_sig00000693
    );
  blk00000003_blk00000536 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000674,
      Q => blk00000003_sig00000692
    );
  blk00000003_blk00000535 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000673,
      Q => blk00000003_sig00000691
    );
  blk00000003_blk00000534 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000672,
      Q => blk00000003_sig00000690
    );
  blk00000003_blk00000533 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000671,
      Q => blk00000003_sig0000068f
    );
  blk00000003_blk00000532 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000670,
      Q => blk00000003_sig0000068e
    );
  blk00000003_blk00000531 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000066f,
      Q => blk00000003_sig0000068d
    );
  blk00000003_blk00000530 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000066e,
      Q => blk00000003_sig0000068c
    );
  blk00000003_blk0000052f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000066d,
      Q => blk00000003_sig0000068b
    );
  blk00000003_blk0000052e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000066c,
      Q => blk00000003_sig0000068a
    );
  blk00000003_blk0000052d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000066b,
      Q => blk00000003_sig00000689
    );
  blk00000003_blk0000052c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000066a,
      Q => blk00000003_sig00000688
    );
  blk00000003_blk0000052b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000669,
      Q => blk00000003_sig00000687
    );
  blk00000003_blk0000052a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000668,
      Q => blk00000003_sig00000686
    );
  blk00000003_blk00000529 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000667,
      Q => blk00000003_sig00000685
    );
  blk00000003_blk00000528 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000666,
      Q => blk00000003_sig00000684
    );
  blk00000003_blk00000527 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000665,
      Q => blk00000003_sig000002fc
    );
  blk00000003_blk00000526 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002c5,
      Q => blk00000003_sig00000683
    );
  blk00000003_blk00000525 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000664,
      Q => blk00000003_sig00000682
    );
  blk00000003_blk00000524 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000663,
      Q => blk00000003_sig00000681
    );
  blk00000003_blk00000523 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000662,
      Q => blk00000003_sig00000680
    );
  blk00000003_blk00000522 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000661,
      Q => blk00000003_sig0000067f
    );
  blk00000003_blk00000521 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000660,
      Q => blk00000003_sig0000067e
    );
  blk00000003_blk00000520 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000065f,
      Q => blk00000003_sig0000067d
    );
  blk00000003_blk0000051f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000065e,
      Q => blk00000003_sig0000067c
    );
  blk00000003_blk0000051e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000065d,
      Q => blk00000003_sig0000067b
    );
  blk00000003_blk0000051d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000065c,
      Q => blk00000003_sig0000067a
    );
  blk00000003_blk0000051c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000065b,
      Q => blk00000003_sig00000679
    );
  blk00000003_blk0000051b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000065a,
      Q => blk00000003_sig00000678
    );
  blk00000003_blk0000051a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000659,
      Q => blk00000003_sig00000677
    );
  blk00000003_blk00000519 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000658,
      Q => blk00000003_sig00000676
    );
  blk00000003_blk00000518 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000657,
      Q => blk00000003_sig00000675
    );
  blk00000003_blk00000517 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000656,
      Q => blk00000003_sig00000674
    );
  blk00000003_blk00000516 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000655,
      Q => blk00000003_sig00000673
    );
  blk00000003_blk00000515 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000654,
      Q => blk00000003_sig00000672
    );
  blk00000003_blk00000514 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000653,
      Q => blk00000003_sig00000671
    );
  blk00000003_blk00000513 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000652,
      Q => blk00000003_sig00000670
    );
  blk00000003_blk00000512 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000651,
      Q => blk00000003_sig0000066f
    );
  blk00000003_blk00000511 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000650,
      Q => blk00000003_sig0000066e
    );
  blk00000003_blk00000510 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000064f,
      Q => blk00000003_sig0000066d
    );
  blk00000003_blk0000050f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000064e,
      Q => blk00000003_sig0000066c
    );
  blk00000003_blk0000050e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000064d,
      Q => blk00000003_sig0000066b
    );
  blk00000003_blk0000050d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000064c,
      Q => blk00000003_sig0000066a
    );
  blk00000003_blk0000050c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000064b,
      Q => blk00000003_sig00000669
    );
  blk00000003_blk0000050b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000064a,
      Q => blk00000003_sig00000668
    );
  blk00000003_blk0000050a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000649,
      Q => blk00000003_sig00000667
    );
  blk00000003_blk00000509 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000648,
      Q => blk00000003_sig00000666
    );
  blk00000003_blk00000508 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000647,
      Q => blk00000003_sig00000665
    );
  blk00000003_blk00000507 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000646,
      Q => blk00000003_sig000002dd
    );
  blk00000003_blk00000506 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002a6,
      Q => blk00000003_sig00000664
    );
  blk00000003_blk00000505 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000645,
      Q => blk00000003_sig00000663
    );
  blk00000003_blk00000504 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000644,
      Q => blk00000003_sig00000662
    );
  blk00000003_blk00000503 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000643,
      Q => blk00000003_sig00000661
    );
  blk00000003_blk00000502 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000642,
      Q => blk00000003_sig00000660
    );
  blk00000003_blk00000501 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000641,
      Q => blk00000003_sig0000065f
    );
  blk00000003_blk00000500 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000640,
      Q => blk00000003_sig0000065e
    );
  blk00000003_blk000004ff : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000063f,
      Q => blk00000003_sig0000065d
    );
  blk00000003_blk000004fe : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000063e,
      Q => blk00000003_sig0000065c
    );
  blk00000003_blk000004fd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000063d,
      Q => blk00000003_sig0000065b
    );
  blk00000003_blk000004fc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000063c,
      Q => blk00000003_sig0000065a
    );
  blk00000003_blk000004fb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000063b,
      Q => blk00000003_sig00000659
    );
  blk00000003_blk000004fa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000063a,
      Q => blk00000003_sig00000658
    );
  blk00000003_blk000004f9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000639,
      Q => blk00000003_sig00000657
    );
  blk00000003_blk000004f8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000638,
      Q => blk00000003_sig00000656
    );
  blk00000003_blk000004f7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000637,
      Q => blk00000003_sig00000655
    );
  blk00000003_blk000004f6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000636,
      Q => blk00000003_sig00000654
    );
  blk00000003_blk000004f5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000635,
      Q => blk00000003_sig00000653
    );
  blk00000003_blk000004f4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000634,
      Q => blk00000003_sig00000652
    );
  blk00000003_blk000004f3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000633,
      Q => blk00000003_sig00000651
    );
  blk00000003_blk000004f2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000632,
      Q => blk00000003_sig00000650
    );
  blk00000003_blk000004f1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000631,
      Q => blk00000003_sig0000064f
    );
  blk00000003_blk000004f0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000630,
      Q => blk00000003_sig0000064e
    );
  blk00000003_blk000004ef : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000062f,
      Q => blk00000003_sig0000064d
    );
  blk00000003_blk000004ee : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000062e,
      Q => blk00000003_sig0000064c
    );
  blk00000003_blk000004ed : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000062d,
      Q => blk00000003_sig0000064b
    );
  blk00000003_blk000004ec : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000062c,
      Q => blk00000003_sig0000064a
    );
  blk00000003_blk000004eb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000062b,
      Q => blk00000003_sig00000649
    );
  blk00000003_blk000004ea : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000062a,
      Q => blk00000003_sig00000648
    );
  blk00000003_blk000004e9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000629,
      Q => blk00000003_sig00000647
    );
  blk00000003_blk000004e8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000628,
      Q => blk00000003_sig00000646
    );
  blk00000003_blk000004e7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000627,
      Q => blk00000003_sig000002be
    );
  blk00000003_blk000004e6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000287,
      Q => blk00000003_sig00000645
    );
  blk00000003_blk000004e5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000008f,
      Q => blk00000003_sig00000644
    );
  blk00000003_blk000004e4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000090,
      Q => blk00000003_sig00000643
    );
  blk00000003_blk000004e3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000091,
      Q => blk00000003_sig00000642
    );
  blk00000003_blk000004e2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000092,
      Q => blk00000003_sig00000641
    );
  blk00000003_blk000004e1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000093,
      Q => blk00000003_sig00000640
    );
  blk00000003_blk000004e0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000094,
      Q => blk00000003_sig0000063f
    );
  blk00000003_blk000004df : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000095,
      Q => blk00000003_sig0000063e
    );
  blk00000003_blk000004de : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000626,
      Q => blk00000003_sig0000063d
    );
  blk00000003_blk000004dd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000625,
      Q => blk00000003_sig0000063c
    );
  blk00000003_blk000004dc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000624,
      Q => blk00000003_sig0000063b
    );
  blk00000003_blk000004db : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000623,
      Q => blk00000003_sig0000063a
    );
  blk00000003_blk000004da : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000622,
      Q => blk00000003_sig00000639
    );
  blk00000003_blk000004d9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000621,
      Q => blk00000003_sig00000638
    );
  blk00000003_blk000004d8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000620,
      Q => blk00000003_sig00000637
    );
  blk00000003_blk000004d7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000061f,
      Q => blk00000003_sig00000636
    );
  blk00000003_blk000004d6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000061e,
      Q => blk00000003_sig00000635
    );
  blk00000003_blk000004d5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000061d,
      Q => blk00000003_sig00000634
    );
  blk00000003_blk000004d4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000061c,
      Q => blk00000003_sig00000633
    );
  blk00000003_blk000004d3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000061b,
      Q => blk00000003_sig00000632
    );
  blk00000003_blk000004d2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000061a,
      Q => blk00000003_sig00000631
    );
  blk00000003_blk000004d1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000619,
      Q => blk00000003_sig00000630
    );
  blk00000003_blk000004d0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000618,
      Q => blk00000003_sig0000062f
    );
  blk00000003_blk000004cf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000617,
      Q => blk00000003_sig0000062e
    );
  blk00000003_blk000004ce : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000616,
      Q => blk00000003_sig0000062d
    );
  blk00000003_blk000004cd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000615,
      Q => blk00000003_sig0000062c
    );
  blk00000003_blk000004cc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000614,
      Q => blk00000003_sig0000062b
    );
  blk00000003_blk000004cb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000613,
      Q => blk00000003_sig0000062a
    );
  blk00000003_blk000004ca : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000612,
      Q => blk00000003_sig00000629
    );
  blk00000003_blk000004c9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000611,
      Q => blk00000003_sig00000628
    );
  blk00000003_blk000004c8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000610,
      Q => blk00000003_sig00000627
    );
  blk00000003_blk000004c7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000060f,
      Q => blk00000003_sig0000029f
    );
  blk00000003_blk000004c6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000060e,
      Q => blk00000003_sig00000626
    );
  blk00000003_blk000004c5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000060d,
      Q => blk00000003_sig00000625
    );
  blk00000003_blk000004c4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000060c,
      Q => blk00000003_sig00000624
    );
  blk00000003_blk000004c3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000060b,
      Q => blk00000003_sig00000623
    );
  blk00000003_blk000004c2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000060a,
      Q => blk00000003_sig00000622
    );
  blk00000003_blk000004c1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000609,
      Q => blk00000003_sig00000621
    );
  blk00000003_blk000004c0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000608,
      Q => blk00000003_sig00000620
    );
  blk00000003_blk000004bf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000607,
      Q => blk00000003_sig0000061f
    );
  blk00000003_blk000004be : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000606,
      Q => blk00000003_sig0000061e
    );
  blk00000003_blk000004bd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000605,
      Q => blk00000003_sig0000061d
    );
  blk00000003_blk000004bc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000604,
      Q => blk00000003_sig0000061c
    );
  blk00000003_blk000004bb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000603,
      Q => blk00000003_sig0000061b
    );
  blk00000003_blk000004ba : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000602,
      Q => blk00000003_sig0000061a
    );
  blk00000003_blk000004b9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000601,
      Q => blk00000003_sig00000619
    );
  blk00000003_blk000004b8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000600,
      Q => blk00000003_sig00000618
    );
  blk00000003_blk000004b7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005ff,
      Q => blk00000003_sig00000617
    );
  blk00000003_blk000004b6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005fe,
      Q => blk00000003_sig00000616
    );
  blk00000003_blk000004b5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005fd,
      Q => blk00000003_sig00000615
    );
  blk00000003_blk000004b4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005fc,
      Q => blk00000003_sig00000614
    );
  blk00000003_blk000004b3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005fb,
      Q => blk00000003_sig00000613
    );
  blk00000003_blk000004b2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005fa,
      Q => blk00000003_sig00000612
    );
  blk00000003_blk000004b1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005f9,
      Q => blk00000003_sig00000611
    );
  blk00000003_blk000004b0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005f8,
      Q => blk00000003_sig00000610
    );
  blk00000003_blk000004af : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005f7,
      Q => blk00000003_sig0000060f
    );
  blk00000003_blk000004ae : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005f6,
      Q => blk00000003_sig00000280
    );
  blk00000003_blk000004ad : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005f5,
      Q => blk00000003_sig0000060e
    );
  blk00000003_blk000004ac : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005f4,
      Q => blk00000003_sig0000060d
    );
  blk00000003_blk000004ab : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005f3,
      Q => blk00000003_sig0000060c
    );
  blk00000003_blk000004aa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005f2,
      Q => blk00000003_sig0000060b
    );
  blk00000003_blk000004a9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005f1,
      Q => blk00000003_sig0000060a
    );
  blk00000003_blk000004a8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005f0,
      Q => blk00000003_sig00000609
    );
  blk00000003_blk000004a7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005ef,
      Q => blk00000003_sig00000608
    );
  blk00000003_blk000004a6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005ee,
      Q => blk00000003_sig00000607
    );
  blk00000003_blk000004a5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005ed,
      Q => blk00000003_sig00000606
    );
  blk00000003_blk000004a4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005ec,
      Q => blk00000003_sig00000605
    );
  blk00000003_blk000004a3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005eb,
      Q => blk00000003_sig00000604
    );
  blk00000003_blk000004a2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005ea,
      Q => blk00000003_sig00000603
    );
  blk00000003_blk000004a1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005e9,
      Q => blk00000003_sig00000602
    );
  blk00000003_blk000004a0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005e8,
      Q => blk00000003_sig00000601
    );
  blk00000003_blk0000049f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005e7,
      Q => blk00000003_sig00000600
    );
  blk00000003_blk0000049e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005e6,
      Q => blk00000003_sig000005ff
    );
  blk00000003_blk0000049d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005e5,
      Q => blk00000003_sig000005fe
    );
  blk00000003_blk0000049c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005e4,
      Q => blk00000003_sig000005fd
    );
  blk00000003_blk0000049b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005e3,
      Q => blk00000003_sig000005fc
    );
  blk00000003_blk0000049a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005e2,
      Q => blk00000003_sig000005fb
    );
  blk00000003_blk00000499 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005e1,
      Q => blk00000003_sig000005fa
    );
  blk00000003_blk00000498 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005e0,
      Q => blk00000003_sig000005f9
    );
  blk00000003_blk00000497 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005df,
      Q => blk00000003_sig000005f8
    );
  blk00000003_blk00000496 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005de,
      Q => blk00000003_sig000005f7
    );
  blk00000003_blk00000495 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005dd,
      Q => blk00000003_sig000005f6
    );
  blk00000003_blk00000494 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005dc,
      Q => blk00000003_sig00000262
    );
  blk00000003_blk00000493 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005db,
      Q => blk00000003_sig000005f5
    );
  blk00000003_blk00000492 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005da,
      Q => blk00000003_sig000005f4
    );
  blk00000003_blk00000491 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005d9,
      Q => blk00000003_sig000005f3
    );
  blk00000003_blk00000490 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005d8,
      Q => blk00000003_sig000005f2
    );
  blk00000003_blk0000048f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005d7,
      Q => blk00000003_sig000005f1
    );
  blk00000003_blk0000048e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005d6,
      Q => blk00000003_sig000005f0
    );
  blk00000003_blk0000048d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005d5,
      Q => blk00000003_sig000005ef
    );
  blk00000003_blk0000048c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005d4,
      Q => blk00000003_sig000005ee
    );
  blk00000003_blk0000048b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005d3,
      Q => blk00000003_sig000005ed
    );
  blk00000003_blk0000048a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005d2,
      Q => blk00000003_sig000005ec
    );
  blk00000003_blk00000489 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005d1,
      Q => blk00000003_sig000005eb
    );
  blk00000003_blk00000488 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005d0,
      Q => blk00000003_sig000005ea
    );
  blk00000003_blk00000487 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005cf,
      Q => blk00000003_sig000005e9
    );
  blk00000003_blk00000486 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005ce,
      Q => blk00000003_sig000005e8
    );
  blk00000003_blk00000485 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005cd,
      Q => blk00000003_sig000005e7
    );
  blk00000003_blk00000484 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005cc,
      Q => blk00000003_sig000005e6
    );
  blk00000003_blk00000483 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005cb,
      Q => blk00000003_sig000005e5
    );
  blk00000003_blk00000482 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005ca,
      Q => blk00000003_sig000005e4
    );
  blk00000003_blk00000481 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005c9,
      Q => blk00000003_sig000005e3
    );
  blk00000003_blk00000480 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005c8,
      Q => blk00000003_sig000005e2
    );
  blk00000003_blk0000047f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005c7,
      Q => blk00000003_sig000005e1
    );
  blk00000003_blk0000047e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005c6,
      Q => blk00000003_sig000005e0
    );
  blk00000003_blk0000047d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005c5,
      Q => blk00000003_sig000005df
    );
  blk00000003_blk0000047c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005c4,
      Q => blk00000003_sig000005de
    );
  blk00000003_blk0000047b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005c3,
      Q => blk00000003_sig000005dd
    );
  blk00000003_blk0000047a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005c2,
      Q => blk00000003_sig000005dc
    );
  blk00000003_blk00000479 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005c1,
      Q => blk00000003_sig00000244
    );
  blk00000003_blk00000478 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005c0,
      Q => blk00000003_sig000005db
    );
  blk00000003_blk00000477 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005bf,
      Q => blk00000003_sig000005da
    );
  blk00000003_blk00000476 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005be,
      Q => blk00000003_sig000005d9
    );
  blk00000003_blk00000475 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005bd,
      Q => blk00000003_sig000005d8
    );
  blk00000003_blk00000474 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005bc,
      Q => blk00000003_sig000005d7
    );
  blk00000003_blk00000473 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005bb,
      Q => blk00000003_sig000005d6
    );
  blk00000003_blk00000472 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005ba,
      Q => blk00000003_sig000005d5
    );
  blk00000003_blk00000471 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005b9,
      Q => blk00000003_sig000005d4
    );
  blk00000003_blk00000470 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005b8,
      Q => blk00000003_sig000005d3
    );
  blk00000003_blk0000046f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005b7,
      Q => blk00000003_sig000005d2
    );
  blk00000003_blk0000046e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005b6,
      Q => blk00000003_sig000005d1
    );
  blk00000003_blk0000046d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005b5,
      Q => blk00000003_sig000005d0
    );
  blk00000003_blk0000046c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005b4,
      Q => blk00000003_sig000005cf
    );
  blk00000003_blk0000046b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005b3,
      Q => blk00000003_sig000005ce
    );
  blk00000003_blk0000046a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005b2,
      Q => blk00000003_sig000005cd
    );
  blk00000003_blk00000469 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005b1,
      Q => blk00000003_sig000005cc
    );
  blk00000003_blk00000468 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005b0,
      Q => blk00000003_sig000005cb
    );
  blk00000003_blk00000467 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005af,
      Q => blk00000003_sig000005ca
    );
  blk00000003_blk00000466 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005ae,
      Q => blk00000003_sig000005c9
    );
  blk00000003_blk00000465 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005ad,
      Q => blk00000003_sig000005c8
    );
  blk00000003_blk00000464 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005ac,
      Q => blk00000003_sig000005c7
    );
  blk00000003_blk00000463 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005ab,
      Q => blk00000003_sig000005c6
    );
  blk00000003_blk00000462 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005aa,
      Q => blk00000003_sig000005c5
    );
  blk00000003_blk00000461 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005a9,
      Q => blk00000003_sig000005c4
    );
  blk00000003_blk00000460 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005a8,
      Q => blk00000003_sig000005c3
    );
  blk00000003_blk0000045f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005a7,
      Q => blk00000003_sig000005c2
    );
  blk00000003_blk0000045e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005a6,
      Q => blk00000003_sig000005c1
    );
  blk00000003_blk0000045d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005a5,
      Q => blk00000003_sig00000226
    );
  blk00000003_blk0000045c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005a4,
      Q => blk00000003_sig000005c0
    );
  blk00000003_blk0000045b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005a3,
      Q => blk00000003_sig000005bf
    );
  blk00000003_blk0000045a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005a2,
      Q => blk00000003_sig000005be
    );
  blk00000003_blk00000459 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005a1,
      Q => blk00000003_sig000005bd
    );
  blk00000003_blk00000458 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000005a0,
      Q => blk00000003_sig000005bc
    );
  blk00000003_blk00000457 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000059f,
      Q => blk00000003_sig000005bb
    );
  blk00000003_blk00000456 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000059e,
      Q => blk00000003_sig000005ba
    );
  blk00000003_blk00000455 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000059d,
      Q => blk00000003_sig000005b9
    );
  blk00000003_blk00000454 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000059c,
      Q => blk00000003_sig000005b8
    );
  blk00000003_blk00000453 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000059b,
      Q => blk00000003_sig000005b7
    );
  blk00000003_blk00000452 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000059a,
      Q => blk00000003_sig000005b6
    );
  blk00000003_blk00000451 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000599,
      Q => blk00000003_sig000005b5
    );
  blk00000003_blk00000450 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000598,
      Q => blk00000003_sig000005b4
    );
  blk00000003_blk0000044f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000597,
      Q => blk00000003_sig000005b3
    );
  blk00000003_blk0000044e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000596,
      Q => blk00000003_sig000005b2
    );
  blk00000003_blk0000044d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000595,
      Q => blk00000003_sig000005b1
    );
  blk00000003_blk0000044c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000594,
      Q => blk00000003_sig000005b0
    );
  blk00000003_blk0000044b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000593,
      Q => blk00000003_sig000005af
    );
  blk00000003_blk0000044a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000592,
      Q => blk00000003_sig000005ae
    );
  blk00000003_blk00000449 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000591,
      Q => blk00000003_sig000005ad
    );
  blk00000003_blk00000448 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000590,
      Q => blk00000003_sig000005ac
    );
  blk00000003_blk00000447 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000058f,
      Q => blk00000003_sig000005ab
    );
  blk00000003_blk00000446 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000058e,
      Q => blk00000003_sig000005aa
    );
  blk00000003_blk00000445 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000058d,
      Q => blk00000003_sig000005a9
    );
  blk00000003_blk00000444 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000058c,
      Q => blk00000003_sig000005a8
    );
  blk00000003_blk00000443 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000058b,
      Q => blk00000003_sig000005a7
    );
  blk00000003_blk00000442 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000058a,
      Q => blk00000003_sig000005a6
    );
  blk00000003_blk00000441 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000589,
      Q => blk00000003_sig000005a5
    );
  blk00000003_blk00000440 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000588,
      Q => blk00000003_sig00000208
    );
  blk00000003_blk0000043f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000587,
      Q => blk00000003_sig000005a4
    );
  blk00000003_blk0000043e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000586,
      Q => blk00000003_sig000005a3
    );
  blk00000003_blk0000043d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000585,
      Q => blk00000003_sig000005a2
    );
  blk00000003_blk0000043c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000584,
      Q => blk00000003_sig000005a1
    );
  blk00000003_blk0000043b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000583,
      Q => blk00000003_sig000005a0
    );
  blk00000003_blk0000043a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000582,
      Q => blk00000003_sig0000059f
    );
  blk00000003_blk00000439 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000581,
      Q => blk00000003_sig0000059e
    );
  blk00000003_blk00000438 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000580,
      Q => blk00000003_sig0000059d
    );
  blk00000003_blk00000437 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000057f,
      Q => blk00000003_sig0000059c
    );
  blk00000003_blk00000436 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000057e,
      Q => blk00000003_sig0000059b
    );
  blk00000003_blk00000435 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000057d,
      Q => blk00000003_sig0000059a
    );
  blk00000003_blk00000434 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000057c,
      Q => blk00000003_sig00000599
    );
  blk00000003_blk00000433 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000057b,
      Q => blk00000003_sig00000598
    );
  blk00000003_blk00000432 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000057a,
      Q => blk00000003_sig00000597
    );
  blk00000003_blk00000431 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000579,
      Q => blk00000003_sig00000596
    );
  blk00000003_blk00000430 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000578,
      Q => blk00000003_sig00000595
    );
  blk00000003_blk0000042f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000577,
      Q => blk00000003_sig00000594
    );
  blk00000003_blk0000042e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000576,
      Q => blk00000003_sig00000593
    );
  blk00000003_blk0000042d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000575,
      Q => blk00000003_sig00000592
    );
  blk00000003_blk0000042c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000574,
      Q => blk00000003_sig00000591
    );
  blk00000003_blk0000042b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000573,
      Q => blk00000003_sig00000590
    );
  blk00000003_blk0000042a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000572,
      Q => blk00000003_sig0000058f
    );
  blk00000003_blk00000429 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000571,
      Q => blk00000003_sig0000058e
    );
  blk00000003_blk00000428 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000570,
      Q => blk00000003_sig0000058d
    );
  blk00000003_blk00000427 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000056f,
      Q => blk00000003_sig0000058c
    );
  blk00000003_blk00000426 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000056e,
      Q => blk00000003_sig0000058b
    );
  blk00000003_blk00000425 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000056d,
      Q => blk00000003_sig0000058a
    );
  blk00000003_blk00000424 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000056c,
      Q => blk00000003_sig00000589
    );
  blk00000003_blk00000423 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000056b,
      Q => blk00000003_sig00000588
    );
  blk00000003_blk00000422 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000056a,
      Q => blk00000003_sig000001ea
    );
  blk00000003_blk00000421 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000019c,
      Q => blk00000003_sig00000587
    );
  blk00000003_blk00000420 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000019b,
      Q => blk00000003_sig00000586
    );
  blk00000003_blk0000041f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000019a,
      Q => blk00000003_sig00000585
    );
  blk00000003_blk0000041e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000199,
      Q => blk00000003_sig00000584
    );
  blk00000003_blk0000041d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000198,
      Q => blk00000003_sig00000583
    );
  blk00000003_blk0000041c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000197,
      Q => blk00000003_sig00000582
    );
  blk00000003_blk0000041b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000196,
      Q => blk00000003_sig00000581
    );
  blk00000003_blk0000041a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000195,
      Q => blk00000003_sig00000580
    );
  blk00000003_blk00000419 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000194,
      Q => blk00000003_sig0000057f
    );
  blk00000003_blk00000418 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000193,
      Q => blk00000003_sig0000057e
    );
  blk00000003_blk00000417 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000192,
      Q => blk00000003_sig0000057d
    );
  blk00000003_blk00000416 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000191,
      Q => blk00000003_sig0000057c
    );
  blk00000003_blk00000415 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000190,
      Q => blk00000003_sig0000057b
    );
  blk00000003_blk00000414 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000018f,
      Q => blk00000003_sig0000057a
    );
  blk00000003_blk00000413 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000018e,
      Q => blk00000003_sig00000579
    );
  blk00000003_blk00000412 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000018d,
      Q => blk00000003_sig00000578
    );
  blk00000003_blk00000411 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000018c,
      Q => blk00000003_sig00000577
    );
  blk00000003_blk00000410 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000018b,
      Q => blk00000003_sig00000576
    );
  blk00000003_blk0000040f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000018a,
      Q => blk00000003_sig00000575
    );
  blk00000003_blk0000040e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000189,
      Q => blk00000003_sig00000574
    );
  blk00000003_blk0000040d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000188,
      Q => blk00000003_sig00000573
    );
  blk00000003_blk0000040c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000187,
      Q => blk00000003_sig00000572
    );
  blk00000003_blk0000040b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000186,
      Q => blk00000003_sig00000571
    );
  blk00000003_blk0000040a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000185,
      Q => blk00000003_sig00000570
    );
  blk00000003_blk00000409 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000184,
      Q => blk00000003_sig0000056f
    );
  blk00000003_blk00000408 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000183,
      Q => blk00000003_sig0000056e
    );
  blk00000003_blk00000407 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000182,
      Q => blk00000003_sig0000056d
    );
  blk00000003_blk00000406 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000181,
      Q => blk00000003_sig0000056c
    );
  blk00000003_blk00000405 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000180,
      Q => blk00000003_sig0000056b
    );
  blk00000003_blk00000404 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000017f,
      Q => blk00000003_sig0000056a
    );
  blk00000003_blk00000403 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000017e,
      Q => blk00000003_sig000001cc
    );
  blk00000003_blk00000402 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000055e,
      Q => blk00000003_sig00000569
    );
  blk00000003_blk00000401 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000054e,
      Q => blk00000003_sig00000568
    );
  blk00000003_blk00000400 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000551,
      Q => blk00000003_sig00000567
    );
  blk00000003_blk000003ff : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000554,
      Q => blk00000003_sig00000566
    );
  blk00000003_blk000003fe : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000557,
      Q => blk00000003_sig00000565
    );
  blk00000003_blk000003fd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000055a,
      Q => blk00000003_sig00000564
    );
  blk00000003_blk000003fc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000055d,
      Q => blk00000003_sig00000563
    );
  blk00000003_blk000003fb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000561,
      Q => blk00000003_sig00000562
    );
  blk00000003_blk000003fa : MUXCY
    port map (
      CI => blk00000003_sig0000055f,
      DI => blk00000003_sig00000096,
      S => blk00000003_sig00000560,
      O => blk00000003_sig0000055b
    );
  blk00000003_blk000003f9 : XORCY
    port map (
      CI => blk00000003_sig0000055f,
      LI => blk00000003_sig00000560,
      O => blk00000003_sig00000561
    );
  blk00000003_blk000003f8 : MUXCY
    port map (
      CI => blk00000003_sig0000054c,
      DI => blk00000003_sig00000549,
      S => blk00000003_sig0000054d,
      O => blk00000003_sig0000055e
    );
  blk00000003_blk000003f7 : MUXCY
    port map (
      CI => blk00000003_sig0000055b,
      DI => blk00000003_sig00000544,
      S => blk00000003_sig0000055c,
      O => blk00000003_sig00000558
    );
  blk00000003_blk000003f6 : MUXCY
    port map (
      CI => blk00000003_sig00000558,
      DI => blk00000003_sig00000545,
      S => blk00000003_sig00000559,
      O => blk00000003_sig00000555
    );
  blk00000003_blk000003f5 : MUXCY
    port map (
      CI => blk00000003_sig00000555,
      DI => blk00000003_sig00000546,
      S => blk00000003_sig00000556,
      O => blk00000003_sig00000552
    );
  blk00000003_blk000003f4 : MUXCY
    port map (
      CI => blk00000003_sig00000552,
      DI => blk00000003_sig00000547,
      S => blk00000003_sig00000553,
      O => blk00000003_sig0000054f
    );
  blk00000003_blk000003f3 : MUXCY
    port map (
      CI => blk00000003_sig0000054f,
      DI => blk00000003_sig00000548,
      S => blk00000003_sig00000550,
      O => blk00000003_sig0000054c
    );
  blk00000003_blk000003f2 : XORCY
    port map (
      CI => blk00000003_sig0000055b,
      LI => blk00000003_sig0000055c,
      O => blk00000003_sig0000055d
    );
  blk00000003_blk000003f1 : XORCY
    port map (
      CI => blk00000003_sig00000558,
      LI => blk00000003_sig00000559,
      O => blk00000003_sig0000055a
    );
  blk00000003_blk000003f0 : XORCY
    port map (
      CI => blk00000003_sig00000555,
      LI => blk00000003_sig00000556,
      O => blk00000003_sig00000557
    );
  blk00000003_blk000003ef : XORCY
    port map (
      CI => blk00000003_sig00000552,
      LI => blk00000003_sig00000553,
      O => blk00000003_sig00000554
    );
  blk00000003_blk000003ee : XORCY
    port map (
      CI => blk00000003_sig0000054f,
      LI => blk00000003_sig00000550,
      O => blk00000003_sig00000551
    );
  blk00000003_blk000003ed : XORCY
    port map (
      CI => blk00000003_sig0000054c,
      LI => blk00000003_sig0000054d,
      O => blk00000003_sig0000054e
    );
  blk00000003_blk000003ec : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000540,
      Q => blk00000003_sig0000054b
    );
  blk00000003_blk000003eb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000530,
      Q => blk00000003_sig0000054a
    );
  blk00000003_blk000003ea : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000533,
      Q => blk00000003_sig00000549
    );
  blk00000003_blk000003e9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000536,
      Q => blk00000003_sig00000548
    );
  blk00000003_blk000003e8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000539,
      Q => blk00000003_sig00000547
    );
  blk00000003_blk000003e7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000053c,
      Q => blk00000003_sig00000546
    );
  blk00000003_blk000003e6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000053f,
      Q => blk00000003_sig00000545
    );
  blk00000003_blk000003e5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000543,
      Q => blk00000003_sig00000544
    );
  blk00000003_blk000003e4 : MUXCY
    port map (
      CI => blk00000003_sig00000541,
      DI => blk00000003_sig00000054,
      S => blk00000003_sig00000542,
      O => blk00000003_sig0000053d
    );
  blk00000003_blk000003e3 : XORCY
    port map (
      CI => blk00000003_sig00000541,
      LI => blk00000003_sig00000542,
      O => blk00000003_sig00000543
    );
  blk00000003_blk000003e2 : MUXCY
    port map (
      CI => blk00000003_sig0000052e,
      DI => blk00000003_sig0000052b,
      S => blk00000003_sig0000052f,
      O => blk00000003_sig00000540
    );
  blk00000003_blk000003e1 : MUXCY
    port map (
      CI => blk00000003_sig0000053d,
      DI => blk00000003_sig00000526,
      S => blk00000003_sig0000053e,
      O => blk00000003_sig0000053a
    );
  blk00000003_blk000003e0 : MUXCY
    port map (
      CI => blk00000003_sig0000053a,
      DI => blk00000003_sig00000527,
      S => blk00000003_sig0000053b,
      O => blk00000003_sig00000537
    );
  blk00000003_blk000003df : MUXCY
    port map (
      CI => blk00000003_sig00000537,
      DI => blk00000003_sig00000528,
      S => blk00000003_sig00000538,
      O => blk00000003_sig00000534
    );
  blk00000003_blk000003de : MUXCY
    port map (
      CI => blk00000003_sig00000534,
      DI => blk00000003_sig00000529,
      S => blk00000003_sig00000535,
      O => blk00000003_sig00000531
    );
  blk00000003_blk000003dd : MUXCY
    port map (
      CI => blk00000003_sig00000531,
      DI => blk00000003_sig0000052a,
      S => blk00000003_sig00000532,
      O => blk00000003_sig0000052e
    );
  blk00000003_blk000003dc : XORCY
    port map (
      CI => blk00000003_sig0000053d,
      LI => blk00000003_sig0000053e,
      O => blk00000003_sig0000053f
    );
  blk00000003_blk000003db : XORCY
    port map (
      CI => blk00000003_sig0000053a,
      LI => blk00000003_sig0000053b,
      O => blk00000003_sig0000053c
    );
  blk00000003_blk000003da : XORCY
    port map (
      CI => blk00000003_sig00000537,
      LI => blk00000003_sig00000538,
      O => blk00000003_sig00000539
    );
  blk00000003_blk000003d9 : XORCY
    port map (
      CI => blk00000003_sig00000534,
      LI => blk00000003_sig00000535,
      O => blk00000003_sig00000536
    );
  blk00000003_blk000003d8 : XORCY
    port map (
      CI => blk00000003_sig00000531,
      LI => blk00000003_sig00000532,
      O => blk00000003_sig00000533
    );
  blk00000003_blk000003d7 : XORCY
    port map (
      CI => blk00000003_sig0000052e,
      LI => blk00000003_sig0000052f,
      O => blk00000003_sig00000530
    );
  blk00000003_blk000003d6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000522,
      Q => blk00000003_sig0000052d
    );
  blk00000003_blk000003d5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000512,
      Q => blk00000003_sig0000052c
    );
  blk00000003_blk000003d4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000515,
      Q => blk00000003_sig0000052b
    );
  blk00000003_blk000003d3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000518,
      Q => blk00000003_sig0000052a
    );
  blk00000003_blk000003d2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000051b,
      Q => blk00000003_sig00000529
    );
  blk00000003_blk000003d1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000051e,
      Q => blk00000003_sig00000528
    );
  blk00000003_blk000003d0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000521,
      Q => blk00000003_sig00000527
    );
  blk00000003_blk000003cf : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000525,
      Q => blk00000003_sig00000526
    );
  blk00000003_blk000003ce : MUXCY
    port map (
      CI => blk00000003_sig00000523,
      DI => blk00000003_sig00000058,
      S => blk00000003_sig00000524,
      O => blk00000003_sig0000051f
    );
  blk00000003_blk000003cd : XORCY
    port map (
      CI => blk00000003_sig00000523,
      LI => blk00000003_sig00000524,
      O => blk00000003_sig00000525
    );
  blk00000003_blk000003cc : MUXCY
    port map (
      CI => blk00000003_sig00000510,
      DI => blk00000003_sig0000050d,
      S => blk00000003_sig00000511,
      O => blk00000003_sig00000522
    );
  blk00000003_blk000003cb : MUXCY
    port map (
      CI => blk00000003_sig0000051f,
      DI => blk00000003_sig00000508,
      S => blk00000003_sig00000520,
      O => blk00000003_sig0000051c
    );
  blk00000003_blk000003ca : MUXCY
    port map (
      CI => blk00000003_sig0000051c,
      DI => blk00000003_sig00000509,
      S => blk00000003_sig0000051d,
      O => blk00000003_sig00000519
    );
  blk00000003_blk000003c9 : MUXCY
    port map (
      CI => blk00000003_sig00000519,
      DI => blk00000003_sig0000050a,
      S => blk00000003_sig0000051a,
      O => blk00000003_sig00000516
    );
  blk00000003_blk000003c8 : MUXCY
    port map (
      CI => blk00000003_sig00000516,
      DI => blk00000003_sig0000050b,
      S => blk00000003_sig00000517,
      O => blk00000003_sig00000513
    );
  blk00000003_blk000003c7 : MUXCY
    port map (
      CI => blk00000003_sig00000513,
      DI => blk00000003_sig0000050c,
      S => blk00000003_sig00000514,
      O => blk00000003_sig00000510
    );
  blk00000003_blk000003c6 : XORCY
    port map (
      CI => blk00000003_sig0000051f,
      LI => blk00000003_sig00000520,
      O => blk00000003_sig00000521
    );
  blk00000003_blk000003c5 : XORCY
    port map (
      CI => blk00000003_sig0000051c,
      LI => blk00000003_sig0000051d,
      O => blk00000003_sig0000051e
    );
  blk00000003_blk000003c4 : XORCY
    port map (
      CI => blk00000003_sig00000519,
      LI => blk00000003_sig0000051a,
      O => blk00000003_sig0000051b
    );
  blk00000003_blk000003c3 : XORCY
    port map (
      CI => blk00000003_sig00000516,
      LI => blk00000003_sig00000517,
      O => blk00000003_sig00000518
    );
  blk00000003_blk000003c2 : XORCY
    port map (
      CI => blk00000003_sig00000513,
      LI => blk00000003_sig00000514,
      O => blk00000003_sig00000515
    );
  blk00000003_blk000003c1 : XORCY
    port map (
      CI => blk00000003_sig00000510,
      LI => blk00000003_sig00000511,
      O => blk00000003_sig00000512
    );
  blk00000003_blk000003c0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000504,
      Q => blk00000003_sig0000050f
    );
  blk00000003_blk000003bf : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004f4,
      Q => blk00000003_sig0000050e
    );
  blk00000003_blk000003be : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004f7,
      Q => blk00000003_sig0000050d
    );
  blk00000003_blk000003bd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004fa,
      Q => blk00000003_sig0000050c
    );
  blk00000003_blk000003bc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004fd,
      Q => blk00000003_sig0000050b
    );
  blk00000003_blk000003bb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000500,
      Q => blk00000003_sig0000050a
    );
  blk00000003_blk000003ba : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000503,
      Q => blk00000003_sig00000509
    );
  blk00000003_blk000003b9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000507,
      Q => blk00000003_sig00000508
    );
  blk00000003_blk000003b8 : MUXCY
    port map (
      CI => blk00000003_sig00000505,
      DI => blk00000003_sig0000005d,
      S => blk00000003_sig00000506,
      O => blk00000003_sig00000501
    );
  blk00000003_blk000003b7 : XORCY
    port map (
      CI => blk00000003_sig00000505,
      LI => blk00000003_sig00000506,
      O => blk00000003_sig00000507
    );
  blk00000003_blk000003b6 : MUXCY
    port map (
      CI => blk00000003_sig000004f2,
      DI => blk00000003_sig000004ef,
      S => blk00000003_sig000004f3,
      O => blk00000003_sig00000504
    );
  blk00000003_blk000003b5 : MUXCY
    port map (
      CI => blk00000003_sig00000501,
      DI => blk00000003_sig000004ea,
      S => blk00000003_sig00000502,
      O => blk00000003_sig000004fe
    );
  blk00000003_blk000003b4 : MUXCY
    port map (
      CI => blk00000003_sig000004fe,
      DI => blk00000003_sig000004eb,
      S => blk00000003_sig000004ff,
      O => blk00000003_sig000004fb
    );
  blk00000003_blk000003b3 : MUXCY
    port map (
      CI => blk00000003_sig000004fb,
      DI => blk00000003_sig000004ec,
      S => blk00000003_sig000004fc,
      O => blk00000003_sig000004f8
    );
  blk00000003_blk000003b2 : MUXCY
    port map (
      CI => blk00000003_sig000004f8,
      DI => blk00000003_sig000004ed,
      S => blk00000003_sig000004f9,
      O => blk00000003_sig000004f5
    );
  blk00000003_blk000003b1 : MUXCY
    port map (
      CI => blk00000003_sig000004f5,
      DI => blk00000003_sig000004ee,
      S => blk00000003_sig000004f6,
      O => blk00000003_sig000004f2
    );
  blk00000003_blk000003b0 : XORCY
    port map (
      CI => blk00000003_sig00000501,
      LI => blk00000003_sig00000502,
      O => blk00000003_sig00000503
    );
  blk00000003_blk000003af : XORCY
    port map (
      CI => blk00000003_sig000004fe,
      LI => blk00000003_sig000004ff,
      O => blk00000003_sig00000500
    );
  blk00000003_blk000003ae : XORCY
    port map (
      CI => blk00000003_sig000004fb,
      LI => blk00000003_sig000004fc,
      O => blk00000003_sig000004fd
    );
  blk00000003_blk000003ad : XORCY
    port map (
      CI => blk00000003_sig000004f8,
      LI => blk00000003_sig000004f9,
      O => blk00000003_sig000004fa
    );
  blk00000003_blk000003ac : XORCY
    port map (
      CI => blk00000003_sig000004f5,
      LI => blk00000003_sig000004f6,
      O => blk00000003_sig000004f7
    );
  blk00000003_blk000003ab : XORCY
    port map (
      CI => blk00000003_sig000004f2,
      LI => blk00000003_sig000004f3,
      O => blk00000003_sig000004f4
    );
  blk00000003_blk000003aa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004e6,
      Q => blk00000003_sig000004f1
    );
  blk00000003_blk000003a9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004d6,
      Q => blk00000003_sig000004f0
    );
  blk00000003_blk000003a8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004d9,
      Q => blk00000003_sig000004ef
    );
  blk00000003_blk000003a7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004dc,
      Q => blk00000003_sig000004ee
    );
  blk00000003_blk000003a6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004df,
      Q => blk00000003_sig000004ed
    );
  blk00000003_blk000003a5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004e2,
      Q => blk00000003_sig000004ec
    );
  blk00000003_blk000003a4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004e5,
      Q => blk00000003_sig000004eb
    );
  blk00000003_blk000003a3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004e9,
      Q => blk00000003_sig000004ea
    );
  blk00000003_blk000003a2 : MUXCY
    port map (
      CI => blk00000003_sig000004e7,
      DI => blk00000003_sig00000063,
      S => blk00000003_sig000004e8,
      O => blk00000003_sig000004e3
    );
  blk00000003_blk000003a1 : XORCY
    port map (
      CI => blk00000003_sig000004e7,
      LI => blk00000003_sig000004e8,
      O => blk00000003_sig000004e9
    );
  blk00000003_blk000003a0 : MUXCY
    port map (
      CI => blk00000003_sig000004d4,
      DI => blk00000003_sig000004d1,
      S => blk00000003_sig000004d5,
      O => blk00000003_sig000004e6
    );
  blk00000003_blk0000039f : MUXCY
    port map (
      CI => blk00000003_sig000004e3,
      DI => blk00000003_sig000004cc,
      S => blk00000003_sig000004e4,
      O => blk00000003_sig000004e0
    );
  blk00000003_blk0000039e : MUXCY
    port map (
      CI => blk00000003_sig000004e0,
      DI => blk00000003_sig000004cd,
      S => blk00000003_sig000004e1,
      O => blk00000003_sig000004dd
    );
  blk00000003_blk0000039d : MUXCY
    port map (
      CI => blk00000003_sig000004dd,
      DI => blk00000003_sig000004ce,
      S => blk00000003_sig000004de,
      O => blk00000003_sig000004da
    );
  blk00000003_blk0000039c : MUXCY
    port map (
      CI => blk00000003_sig000004da,
      DI => blk00000003_sig000004cf,
      S => blk00000003_sig000004db,
      O => blk00000003_sig000004d7
    );
  blk00000003_blk0000039b : MUXCY
    port map (
      CI => blk00000003_sig000004d7,
      DI => blk00000003_sig000004d0,
      S => blk00000003_sig000004d8,
      O => blk00000003_sig000004d4
    );
  blk00000003_blk0000039a : XORCY
    port map (
      CI => blk00000003_sig000004e3,
      LI => blk00000003_sig000004e4,
      O => blk00000003_sig000004e5
    );
  blk00000003_blk00000399 : XORCY
    port map (
      CI => blk00000003_sig000004e0,
      LI => blk00000003_sig000004e1,
      O => blk00000003_sig000004e2
    );
  blk00000003_blk00000398 : XORCY
    port map (
      CI => blk00000003_sig000004dd,
      LI => blk00000003_sig000004de,
      O => blk00000003_sig000004df
    );
  blk00000003_blk00000397 : XORCY
    port map (
      CI => blk00000003_sig000004da,
      LI => blk00000003_sig000004db,
      O => blk00000003_sig000004dc
    );
  blk00000003_blk00000396 : XORCY
    port map (
      CI => blk00000003_sig000004d7,
      LI => blk00000003_sig000004d8,
      O => blk00000003_sig000004d9
    );
  blk00000003_blk00000395 : XORCY
    port map (
      CI => blk00000003_sig000004d4,
      LI => blk00000003_sig000004d5,
      O => blk00000003_sig000004d6
    );
  blk00000003_blk00000394 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004c8,
      Q => blk00000003_sig000004d3
    );
  blk00000003_blk00000393 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004b8,
      Q => blk00000003_sig000004d2
    );
  blk00000003_blk00000392 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004bb,
      Q => blk00000003_sig000004d1
    );
  blk00000003_blk00000391 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004be,
      Q => blk00000003_sig000004d0
    );
  blk00000003_blk00000390 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004c1,
      Q => blk00000003_sig000004cf
    );
  blk00000003_blk0000038f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004c4,
      Q => blk00000003_sig000004ce
    );
  blk00000003_blk0000038e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004c7,
      Q => blk00000003_sig000004cd
    );
  blk00000003_blk0000038d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004cb,
      Q => blk00000003_sig000004cc
    );
  blk00000003_blk0000038c : MUXCY
    port map (
      CI => blk00000003_sig000004c9,
      DI => blk00000003_sig0000006a,
      S => blk00000003_sig000004ca,
      O => blk00000003_sig000004c5
    );
  blk00000003_blk0000038b : XORCY
    port map (
      CI => blk00000003_sig000004c9,
      LI => blk00000003_sig000004ca,
      O => blk00000003_sig000004cb
    );
  blk00000003_blk0000038a : MUXCY
    port map (
      CI => blk00000003_sig000004b6,
      DI => blk00000003_sig000004b3,
      S => blk00000003_sig000004b7,
      O => blk00000003_sig000004c8
    );
  blk00000003_blk00000389 : MUXCY
    port map (
      CI => blk00000003_sig000004c5,
      DI => blk00000003_sig000004ae,
      S => blk00000003_sig000004c6,
      O => blk00000003_sig000004c2
    );
  blk00000003_blk00000388 : MUXCY
    port map (
      CI => blk00000003_sig000004c2,
      DI => blk00000003_sig000004af,
      S => blk00000003_sig000004c3,
      O => blk00000003_sig000004bf
    );
  blk00000003_blk00000387 : MUXCY
    port map (
      CI => blk00000003_sig000004bf,
      DI => blk00000003_sig000004b0,
      S => blk00000003_sig000004c0,
      O => blk00000003_sig000004bc
    );
  blk00000003_blk00000386 : MUXCY
    port map (
      CI => blk00000003_sig000004bc,
      DI => blk00000003_sig000004b1,
      S => blk00000003_sig000004bd,
      O => blk00000003_sig000004b9
    );
  blk00000003_blk00000385 : MUXCY
    port map (
      CI => blk00000003_sig000004b9,
      DI => blk00000003_sig000004b2,
      S => blk00000003_sig000004ba,
      O => blk00000003_sig000004b6
    );
  blk00000003_blk00000384 : XORCY
    port map (
      CI => blk00000003_sig000004c5,
      LI => blk00000003_sig000004c6,
      O => blk00000003_sig000004c7
    );
  blk00000003_blk00000383 : XORCY
    port map (
      CI => blk00000003_sig000004c2,
      LI => blk00000003_sig000004c3,
      O => blk00000003_sig000004c4
    );
  blk00000003_blk00000382 : XORCY
    port map (
      CI => blk00000003_sig000004bf,
      LI => blk00000003_sig000004c0,
      O => blk00000003_sig000004c1
    );
  blk00000003_blk00000381 : XORCY
    port map (
      CI => blk00000003_sig000004bc,
      LI => blk00000003_sig000004bd,
      O => blk00000003_sig000004be
    );
  blk00000003_blk00000380 : XORCY
    port map (
      CI => blk00000003_sig000004b9,
      LI => blk00000003_sig000004ba,
      O => blk00000003_sig000004bb
    );
  blk00000003_blk0000037f : XORCY
    port map (
      CI => blk00000003_sig000004b6,
      LI => blk00000003_sig000004b7,
      O => blk00000003_sig000004b8
    );
  blk00000003_blk0000037e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004aa,
      Q => blk00000003_sig000004b5
    );
  blk00000003_blk0000037d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000049a,
      Q => blk00000003_sig000004b4
    );
  blk00000003_blk0000037c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000049d,
      Q => blk00000003_sig000004b3
    );
  blk00000003_blk0000037b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004a0,
      Q => blk00000003_sig000004b2
    );
  blk00000003_blk0000037a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004a3,
      Q => blk00000003_sig000004b1
    );
  blk00000003_blk00000379 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004a6,
      Q => blk00000003_sig000004b0
    );
  blk00000003_blk00000378 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004a9,
      Q => blk00000003_sig000004af
    );
  blk00000003_blk00000377 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000004ad,
      Q => blk00000003_sig000004ae
    );
  blk00000003_blk00000376 : MUXCY
    port map (
      CI => blk00000003_sig000004ab,
      DI => blk00000003_sig00000072,
      S => blk00000003_sig000004ac,
      O => blk00000003_sig000004a7
    );
  blk00000003_blk00000375 : XORCY
    port map (
      CI => blk00000003_sig000004ab,
      LI => blk00000003_sig000004ac,
      O => blk00000003_sig000004ad
    );
  blk00000003_blk00000374 : MUXCY
    port map (
      CI => blk00000003_sig00000498,
      DI => blk00000003_sig00000495,
      S => blk00000003_sig00000499,
      O => blk00000003_sig000004aa
    );
  blk00000003_blk00000373 : MUXCY
    port map (
      CI => blk00000003_sig000004a7,
      DI => blk00000003_sig00000490,
      S => blk00000003_sig000004a8,
      O => blk00000003_sig000004a4
    );
  blk00000003_blk00000372 : MUXCY
    port map (
      CI => blk00000003_sig000004a4,
      DI => blk00000003_sig00000491,
      S => blk00000003_sig000004a5,
      O => blk00000003_sig000004a1
    );
  blk00000003_blk00000371 : MUXCY
    port map (
      CI => blk00000003_sig000004a1,
      DI => blk00000003_sig00000492,
      S => blk00000003_sig000004a2,
      O => blk00000003_sig0000049e
    );
  blk00000003_blk00000370 : MUXCY
    port map (
      CI => blk00000003_sig0000049e,
      DI => blk00000003_sig00000493,
      S => blk00000003_sig0000049f,
      O => blk00000003_sig0000049b
    );
  blk00000003_blk0000036f : MUXCY
    port map (
      CI => blk00000003_sig0000049b,
      DI => blk00000003_sig00000494,
      S => blk00000003_sig0000049c,
      O => blk00000003_sig00000498
    );
  blk00000003_blk0000036e : XORCY
    port map (
      CI => blk00000003_sig000004a7,
      LI => blk00000003_sig000004a8,
      O => blk00000003_sig000004a9
    );
  blk00000003_blk0000036d : XORCY
    port map (
      CI => blk00000003_sig000004a4,
      LI => blk00000003_sig000004a5,
      O => blk00000003_sig000004a6
    );
  blk00000003_blk0000036c : XORCY
    port map (
      CI => blk00000003_sig000004a1,
      LI => blk00000003_sig000004a2,
      O => blk00000003_sig000004a3
    );
  blk00000003_blk0000036b : XORCY
    port map (
      CI => blk00000003_sig0000049e,
      LI => blk00000003_sig0000049f,
      O => blk00000003_sig000004a0
    );
  blk00000003_blk0000036a : XORCY
    port map (
      CI => blk00000003_sig0000049b,
      LI => blk00000003_sig0000049c,
      O => blk00000003_sig0000049d
    );
  blk00000003_blk00000369 : XORCY
    port map (
      CI => blk00000003_sig00000498,
      LI => blk00000003_sig00000499,
      O => blk00000003_sig0000049a
    );
  blk00000003_blk00000368 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000048b,
      Q => blk00000003_sig00000497
    );
  blk00000003_blk00000367 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000047b,
      Q => blk00000003_sig00000496
    );
  blk00000003_blk00000366 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000047e,
      Q => blk00000003_sig00000495
    );
  blk00000003_blk00000365 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000481,
      Q => blk00000003_sig00000494
    );
  blk00000003_blk00000364 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000484,
      Q => blk00000003_sig00000493
    );
  blk00000003_blk00000363 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000487,
      Q => blk00000003_sig00000492
    );
  blk00000003_blk00000362 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000048a,
      Q => blk00000003_sig00000491
    );
  blk00000003_blk00000361 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000048e,
      Q => blk00000003_sig00000490
    );
  blk00000003_blk00000360 : MUXCY
    port map (
      CI => blk00000003_sig0000048c,
      DI => blk00000003_sig0000048f,
      S => blk00000003_sig0000048d,
      O => blk00000003_sig00000488
    );
  blk00000003_blk0000035f : XORCY
    port map (
      CI => blk00000003_sig0000048c,
      LI => blk00000003_sig0000048d,
      O => blk00000003_sig0000048e
    );
  blk00000003_blk0000035e : MUXCY
    port map (
      CI => blk00000003_sig00000479,
      DI => blk00000003_sig00000476,
      S => blk00000003_sig0000047a,
      O => blk00000003_sig0000048b
    );
  blk00000003_blk0000035d : MUXCY
    port map (
      CI => blk00000003_sig00000488,
      DI => blk00000003_sig00000471,
      S => blk00000003_sig00000489,
      O => blk00000003_sig00000485
    );
  blk00000003_blk0000035c : MUXCY
    port map (
      CI => blk00000003_sig00000485,
      DI => blk00000003_sig00000472,
      S => blk00000003_sig00000486,
      O => blk00000003_sig00000482
    );
  blk00000003_blk0000035b : MUXCY
    port map (
      CI => blk00000003_sig00000482,
      DI => blk00000003_sig00000473,
      S => blk00000003_sig00000483,
      O => blk00000003_sig0000047f
    );
  blk00000003_blk0000035a : MUXCY
    port map (
      CI => blk00000003_sig0000047f,
      DI => blk00000003_sig00000474,
      S => blk00000003_sig00000480,
      O => blk00000003_sig0000047c
    );
  blk00000003_blk00000359 : MUXCY
    port map (
      CI => blk00000003_sig0000047c,
      DI => blk00000003_sig00000475,
      S => blk00000003_sig0000047d,
      O => blk00000003_sig00000479
    );
  blk00000003_blk00000358 : XORCY
    port map (
      CI => blk00000003_sig00000488,
      LI => blk00000003_sig00000489,
      O => blk00000003_sig0000048a
    );
  blk00000003_blk00000357 : XORCY
    port map (
      CI => blk00000003_sig00000485,
      LI => blk00000003_sig00000486,
      O => blk00000003_sig00000487
    );
  blk00000003_blk00000356 : XORCY
    port map (
      CI => blk00000003_sig00000482,
      LI => blk00000003_sig00000483,
      O => blk00000003_sig00000484
    );
  blk00000003_blk00000355 : XORCY
    port map (
      CI => blk00000003_sig0000047f,
      LI => blk00000003_sig00000480,
      O => blk00000003_sig00000481
    );
  blk00000003_blk00000354 : XORCY
    port map (
      CI => blk00000003_sig0000047c,
      LI => blk00000003_sig0000047d,
      O => blk00000003_sig0000047e
    );
  blk00000003_blk00000353 : XORCY
    port map (
      CI => blk00000003_sig00000479,
      LI => blk00000003_sig0000047a,
      O => blk00000003_sig0000047b
    );
  blk00000003_blk00000352 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000046c,
      Q => blk00000003_sig00000478
    );
  blk00000003_blk00000351 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000045c,
      Q => blk00000003_sig00000477
    );
  blk00000003_blk00000350 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000045f,
      Q => blk00000003_sig00000476
    );
  blk00000003_blk0000034f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000462,
      Q => blk00000003_sig00000475
    );
  blk00000003_blk0000034e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000465,
      Q => blk00000003_sig00000474
    );
  blk00000003_blk0000034d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000468,
      Q => blk00000003_sig00000473
    );
  blk00000003_blk0000034c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000046b,
      Q => blk00000003_sig00000472
    );
  blk00000003_blk0000034b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000046f,
      Q => blk00000003_sig00000471
    );
  blk00000003_blk0000034a : MUXCY
    port map (
      CI => blk00000003_sig0000046d,
      DI => blk00000003_sig00000470,
      S => blk00000003_sig0000046e,
      O => blk00000003_sig00000469
    );
  blk00000003_blk00000349 : XORCY
    port map (
      CI => blk00000003_sig0000046d,
      LI => blk00000003_sig0000046e,
      O => blk00000003_sig0000046f
    );
  blk00000003_blk00000348 : MUXCY
    port map (
      CI => blk00000003_sig0000045a,
      DI => blk00000003_sig00000457,
      S => blk00000003_sig0000045b,
      O => blk00000003_sig0000046c
    );
  blk00000003_blk00000347 : MUXCY
    port map (
      CI => blk00000003_sig00000469,
      DI => blk00000003_sig00000452,
      S => blk00000003_sig0000046a,
      O => blk00000003_sig00000466
    );
  blk00000003_blk00000346 : MUXCY
    port map (
      CI => blk00000003_sig00000466,
      DI => blk00000003_sig00000453,
      S => blk00000003_sig00000467,
      O => blk00000003_sig00000463
    );
  blk00000003_blk00000345 : MUXCY
    port map (
      CI => blk00000003_sig00000463,
      DI => blk00000003_sig00000454,
      S => blk00000003_sig00000464,
      O => blk00000003_sig00000460
    );
  blk00000003_blk00000344 : MUXCY
    port map (
      CI => blk00000003_sig00000460,
      DI => blk00000003_sig00000455,
      S => blk00000003_sig00000461,
      O => blk00000003_sig0000045d
    );
  blk00000003_blk00000343 : MUXCY
    port map (
      CI => blk00000003_sig0000045d,
      DI => blk00000003_sig00000456,
      S => blk00000003_sig0000045e,
      O => blk00000003_sig0000045a
    );
  blk00000003_blk00000342 : XORCY
    port map (
      CI => blk00000003_sig00000469,
      LI => blk00000003_sig0000046a,
      O => blk00000003_sig0000046b
    );
  blk00000003_blk00000341 : XORCY
    port map (
      CI => blk00000003_sig00000466,
      LI => blk00000003_sig00000467,
      O => blk00000003_sig00000468
    );
  blk00000003_blk00000340 : XORCY
    port map (
      CI => blk00000003_sig00000463,
      LI => blk00000003_sig00000464,
      O => blk00000003_sig00000465
    );
  blk00000003_blk0000033f : XORCY
    port map (
      CI => blk00000003_sig00000460,
      LI => blk00000003_sig00000461,
      O => blk00000003_sig00000462
    );
  blk00000003_blk0000033e : XORCY
    port map (
      CI => blk00000003_sig0000045d,
      LI => blk00000003_sig0000045e,
      O => blk00000003_sig0000045f
    );
  blk00000003_blk0000033d : XORCY
    port map (
      CI => blk00000003_sig0000045a,
      LI => blk00000003_sig0000045b,
      O => blk00000003_sig0000045c
    );
  blk00000003_blk0000033c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000044d,
      Q => blk00000003_sig00000459
    );
  blk00000003_blk0000033b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000043d,
      Q => blk00000003_sig00000458
    );
  blk00000003_blk0000033a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000440,
      Q => blk00000003_sig00000457
    );
  blk00000003_blk00000339 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000443,
      Q => blk00000003_sig00000456
    );
  blk00000003_blk00000338 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000446,
      Q => blk00000003_sig00000455
    );
  blk00000003_blk00000337 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000449,
      Q => blk00000003_sig00000454
    );
  blk00000003_blk00000336 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000044c,
      Q => blk00000003_sig00000453
    );
  blk00000003_blk00000335 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000450,
      Q => blk00000003_sig00000452
    );
  blk00000003_blk00000334 : MUXCY
    port map (
      CI => blk00000003_sig0000044e,
      DI => blk00000003_sig00000451,
      S => blk00000003_sig0000044f,
      O => blk00000003_sig0000044a
    );
  blk00000003_blk00000333 : XORCY
    port map (
      CI => blk00000003_sig0000044e,
      LI => blk00000003_sig0000044f,
      O => blk00000003_sig00000450
    );
  blk00000003_blk00000332 : MUXCY
    port map (
      CI => blk00000003_sig0000043b,
      DI => blk00000003_sig00000438,
      S => blk00000003_sig0000043c,
      O => blk00000003_sig0000044d
    );
  blk00000003_blk00000331 : MUXCY
    port map (
      CI => blk00000003_sig0000044a,
      DI => blk00000003_sig00000433,
      S => blk00000003_sig0000044b,
      O => blk00000003_sig00000447
    );
  blk00000003_blk00000330 : MUXCY
    port map (
      CI => blk00000003_sig00000447,
      DI => blk00000003_sig00000434,
      S => blk00000003_sig00000448,
      O => blk00000003_sig00000444
    );
  blk00000003_blk0000032f : MUXCY
    port map (
      CI => blk00000003_sig00000444,
      DI => blk00000003_sig00000435,
      S => blk00000003_sig00000445,
      O => blk00000003_sig00000441
    );
  blk00000003_blk0000032e : MUXCY
    port map (
      CI => blk00000003_sig00000441,
      DI => blk00000003_sig00000436,
      S => blk00000003_sig00000442,
      O => blk00000003_sig0000043e
    );
  blk00000003_blk0000032d : MUXCY
    port map (
      CI => blk00000003_sig0000043e,
      DI => blk00000003_sig00000437,
      S => blk00000003_sig0000043f,
      O => blk00000003_sig0000043b
    );
  blk00000003_blk0000032c : XORCY
    port map (
      CI => blk00000003_sig0000044a,
      LI => blk00000003_sig0000044b,
      O => blk00000003_sig0000044c
    );
  blk00000003_blk0000032b : XORCY
    port map (
      CI => blk00000003_sig00000447,
      LI => blk00000003_sig00000448,
      O => blk00000003_sig00000449
    );
  blk00000003_blk0000032a : XORCY
    port map (
      CI => blk00000003_sig00000444,
      LI => blk00000003_sig00000445,
      O => blk00000003_sig00000446
    );
  blk00000003_blk00000329 : XORCY
    port map (
      CI => blk00000003_sig00000441,
      LI => blk00000003_sig00000442,
      O => blk00000003_sig00000443
    );
  blk00000003_blk00000328 : XORCY
    port map (
      CI => blk00000003_sig0000043e,
      LI => blk00000003_sig0000043f,
      O => blk00000003_sig00000440
    );
  blk00000003_blk00000327 : XORCY
    port map (
      CI => blk00000003_sig0000043b,
      LI => blk00000003_sig0000043c,
      O => blk00000003_sig0000043d
    );
  blk00000003_blk00000326 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000042e,
      Q => blk00000003_sig0000043a
    );
  blk00000003_blk00000325 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000041e,
      Q => blk00000003_sig00000439
    );
  blk00000003_blk00000324 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000421,
      Q => blk00000003_sig00000438
    );
  blk00000003_blk00000323 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000424,
      Q => blk00000003_sig00000437
    );
  blk00000003_blk00000322 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000427,
      Q => blk00000003_sig00000436
    );
  blk00000003_blk00000321 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000042a,
      Q => blk00000003_sig00000435
    );
  blk00000003_blk00000320 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000042d,
      Q => blk00000003_sig00000434
    );
  blk00000003_blk0000031f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000431,
      Q => blk00000003_sig00000433
    );
  blk00000003_blk0000031e : MUXCY
    port map (
      CI => blk00000003_sig0000042f,
      DI => blk00000003_sig00000432,
      S => blk00000003_sig00000430,
      O => blk00000003_sig0000042b
    );
  blk00000003_blk0000031d : XORCY
    port map (
      CI => blk00000003_sig0000042f,
      LI => blk00000003_sig00000430,
      O => blk00000003_sig00000431
    );
  blk00000003_blk0000031c : MUXCY
    port map (
      CI => blk00000003_sig0000041c,
      DI => blk00000003_sig00000419,
      S => blk00000003_sig0000041d,
      O => blk00000003_sig0000042e
    );
  blk00000003_blk0000031b : MUXCY
    port map (
      CI => blk00000003_sig0000042b,
      DI => blk00000003_sig00000414,
      S => blk00000003_sig0000042c,
      O => blk00000003_sig00000428
    );
  blk00000003_blk0000031a : MUXCY
    port map (
      CI => blk00000003_sig00000428,
      DI => blk00000003_sig00000415,
      S => blk00000003_sig00000429,
      O => blk00000003_sig00000425
    );
  blk00000003_blk00000319 : MUXCY
    port map (
      CI => blk00000003_sig00000425,
      DI => blk00000003_sig00000416,
      S => blk00000003_sig00000426,
      O => blk00000003_sig00000422
    );
  blk00000003_blk00000318 : MUXCY
    port map (
      CI => blk00000003_sig00000422,
      DI => blk00000003_sig00000417,
      S => blk00000003_sig00000423,
      O => blk00000003_sig0000041f
    );
  blk00000003_blk00000317 : MUXCY
    port map (
      CI => blk00000003_sig0000041f,
      DI => blk00000003_sig00000418,
      S => blk00000003_sig00000420,
      O => blk00000003_sig0000041c
    );
  blk00000003_blk00000316 : XORCY
    port map (
      CI => blk00000003_sig0000042b,
      LI => blk00000003_sig0000042c,
      O => blk00000003_sig0000042d
    );
  blk00000003_blk00000315 : XORCY
    port map (
      CI => blk00000003_sig00000428,
      LI => blk00000003_sig00000429,
      O => blk00000003_sig0000042a
    );
  blk00000003_blk00000314 : XORCY
    port map (
      CI => blk00000003_sig00000425,
      LI => blk00000003_sig00000426,
      O => blk00000003_sig00000427
    );
  blk00000003_blk00000313 : XORCY
    port map (
      CI => blk00000003_sig00000422,
      LI => blk00000003_sig00000423,
      O => blk00000003_sig00000424
    );
  blk00000003_blk00000312 : XORCY
    port map (
      CI => blk00000003_sig0000041f,
      LI => blk00000003_sig00000420,
      O => blk00000003_sig00000421
    );
  blk00000003_blk00000311 : XORCY
    port map (
      CI => blk00000003_sig0000041c,
      LI => blk00000003_sig0000041d,
      O => blk00000003_sig0000041e
    );
  blk00000003_blk00000310 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000040f,
      Q => blk00000003_sig0000041b
    );
  blk00000003_blk0000030f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003ff,
      Q => blk00000003_sig0000041a
    );
  blk00000003_blk0000030e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000402,
      Q => blk00000003_sig00000419
    );
  blk00000003_blk0000030d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000405,
      Q => blk00000003_sig00000418
    );
  blk00000003_blk0000030c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000408,
      Q => blk00000003_sig00000417
    );
  blk00000003_blk0000030b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000040b,
      Q => blk00000003_sig00000416
    );
  blk00000003_blk0000030a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000040e,
      Q => blk00000003_sig00000415
    );
  blk00000003_blk00000309 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000412,
      Q => blk00000003_sig00000414
    );
  blk00000003_blk00000308 : MUXCY
    port map (
      CI => blk00000003_sig00000410,
      DI => blk00000003_sig00000413,
      S => blk00000003_sig00000411,
      O => blk00000003_sig0000040c
    );
  blk00000003_blk00000307 : XORCY
    port map (
      CI => blk00000003_sig00000410,
      LI => blk00000003_sig00000411,
      O => blk00000003_sig00000412
    );
  blk00000003_blk00000306 : MUXCY
    port map (
      CI => blk00000003_sig000003fd,
      DI => blk00000003_sig000003fa,
      S => blk00000003_sig000003fe,
      O => blk00000003_sig0000040f
    );
  blk00000003_blk00000305 : MUXCY
    port map (
      CI => blk00000003_sig0000040c,
      DI => blk00000003_sig000003f5,
      S => blk00000003_sig0000040d,
      O => blk00000003_sig00000409
    );
  blk00000003_blk00000304 : MUXCY
    port map (
      CI => blk00000003_sig00000409,
      DI => blk00000003_sig000003f6,
      S => blk00000003_sig0000040a,
      O => blk00000003_sig00000406
    );
  blk00000003_blk00000303 : MUXCY
    port map (
      CI => blk00000003_sig00000406,
      DI => blk00000003_sig000003f7,
      S => blk00000003_sig00000407,
      O => blk00000003_sig00000403
    );
  blk00000003_blk00000302 : MUXCY
    port map (
      CI => blk00000003_sig00000403,
      DI => blk00000003_sig000003f8,
      S => blk00000003_sig00000404,
      O => blk00000003_sig00000400
    );
  blk00000003_blk00000301 : MUXCY
    port map (
      CI => blk00000003_sig00000400,
      DI => blk00000003_sig000003f9,
      S => blk00000003_sig00000401,
      O => blk00000003_sig000003fd
    );
  blk00000003_blk00000300 : XORCY
    port map (
      CI => blk00000003_sig0000040c,
      LI => blk00000003_sig0000040d,
      O => blk00000003_sig0000040e
    );
  blk00000003_blk000002ff : XORCY
    port map (
      CI => blk00000003_sig00000409,
      LI => blk00000003_sig0000040a,
      O => blk00000003_sig0000040b
    );
  blk00000003_blk000002fe : XORCY
    port map (
      CI => blk00000003_sig00000406,
      LI => blk00000003_sig00000407,
      O => blk00000003_sig00000408
    );
  blk00000003_blk000002fd : XORCY
    port map (
      CI => blk00000003_sig00000403,
      LI => blk00000003_sig00000404,
      O => blk00000003_sig00000405
    );
  blk00000003_blk000002fc : XORCY
    port map (
      CI => blk00000003_sig00000400,
      LI => blk00000003_sig00000401,
      O => blk00000003_sig00000402
    );
  blk00000003_blk000002fb : XORCY
    port map (
      CI => blk00000003_sig000003fd,
      LI => blk00000003_sig000003fe,
      O => blk00000003_sig000003ff
    );
  blk00000003_blk000002fa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003f0,
      Q => blk00000003_sig000003fc
    );
  blk00000003_blk000002f9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003e0,
      Q => blk00000003_sig000003fb
    );
  blk00000003_blk000002f8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003e3,
      Q => blk00000003_sig000003fa
    );
  blk00000003_blk000002f7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003e6,
      Q => blk00000003_sig000003f9
    );
  blk00000003_blk000002f6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003e9,
      Q => blk00000003_sig000003f8
    );
  blk00000003_blk000002f5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003ec,
      Q => blk00000003_sig000003f7
    );
  blk00000003_blk000002f4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003ef,
      Q => blk00000003_sig000003f6
    );
  blk00000003_blk000002f3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003f3,
      Q => blk00000003_sig000003f5
    );
  blk00000003_blk000002f2 : MUXCY
    port map (
      CI => blk00000003_sig000003f1,
      DI => blk00000003_sig000003f4,
      S => blk00000003_sig000003f2,
      O => blk00000003_sig000003ed
    );
  blk00000003_blk000002f1 : XORCY
    port map (
      CI => blk00000003_sig000003f1,
      LI => blk00000003_sig000003f2,
      O => blk00000003_sig000003f3
    );
  blk00000003_blk000002f0 : MUXCY
    port map (
      CI => blk00000003_sig000003de,
      DI => blk00000003_sig000003db,
      S => blk00000003_sig000003df,
      O => blk00000003_sig000003f0
    );
  blk00000003_blk000002ef : MUXCY
    port map (
      CI => blk00000003_sig000003ed,
      DI => blk00000003_sig000003d6,
      S => blk00000003_sig000003ee,
      O => blk00000003_sig000003ea
    );
  blk00000003_blk000002ee : MUXCY
    port map (
      CI => blk00000003_sig000003ea,
      DI => blk00000003_sig000003d7,
      S => blk00000003_sig000003eb,
      O => blk00000003_sig000003e7
    );
  blk00000003_blk000002ed : MUXCY
    port map (
      CI => blk00000003_sig000003e7,
      DI => blk00000003_sig000003d8,
      S => blk00000003_sig000003e8,
      O => blk00000003_sig000003e4
    );
  blk00000003_blk000002ec : MUXCY
    port map (
      CI => blk00000003_sig000003e4,
      DI => blk00000003_sig000003d9,
      S => blk00000003_sig000003e5,
      O => blk00000003_sig000003e1
    );
  blk00000003_blk000002eb : MUXCY
    port map (
      CI => blk00000003_sig000003e1,
      DI => blk00000003_sig000003da,
      S => blk00000003_sig000003e2,
      O => blk00000003_sig000003de
    );
  blk00000003_blk000002ea : XORCY
    port map (
      CI => blk00000003_sig000003ed,
      LI => blk00000003_sig000003ee,
      O => blk00000003_sig000003ef
    );
  blk00000003_blk000002e9 : XORCY
    port map (
      CI => blk00000003_sig000003ea,
      LI => blk00000003_sig000003eb,
      O => blk00000003_sig000003ec
    );
  blk00000003_blk000002e8 : XORCY
    port map (
      CI => blk00000003_sig000003e7,
      LI => blk00000003_sig000003e8,
      O => blk00000003_sig000003e9
    );
  blk00000003_blk000002e7 : XORCY
    port map (
      CI => blk00000003_sig000003e4,
      LI => blk00000003_sig000003e5,
      O => blk00000003_sig000003e6
    );
  blk00000003_blk000002e6 : XORCY
    port map (
      CI => blk00000003_sig000003e1,
      LI => blk00000003_sig000003e2,
      O => blk00000003_sig000003e3
    );
  blk00000003_blk000002e5 : XORCY
    port map (
      CI => blk00000003_sig000003de,
      LI => blk00000003_sig000003df,
      O => blk00000003_sig000003e0
    );
  blk00000003_blk000002e4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003d1,
      Q => blk00000003_sig000003dd
    );
  blk00000003_blk000002e3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003c1,
      Q => blk00000003_sig000003dc
    );
  blk00000003_blk000002e2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003c4,
      Q => blk00000003_sig000003db
    );
  blk00000003_blk000002e1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003c7,
      Q => blk00000003_sig000003da
    );
  blk00000003_blk000002e0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003ca,
      Q => blk00000003_sig000003d9
    );
  blk00000003_blk000002df : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003cd,
      Q => blk00000003_sig000003d8
    );
  blk00000003_blk000002de : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003d0,
      Q => blk00000003_sig000003d7
    );
  blk00000003_blk000002dd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003d4,
      Q => blk00000003_sig000003d6
    );
  blk00000003_blk000002dc : MUXCY
    port map (
      CI => blk00000003_sig000003d2,
      DI => blk00000003_sig000003d5,
      S => blk00000003_sig000003d3,
      O => blk00000003_sig000003ce
    );
  blk00000003_blk000002db : XORCY
    port map (
      CI => blk00000003_sig000003d2,
      LI => blk00000003_sig000003d3,
      O => blk00000003_sig000003d4
    );
  blk00000003_blk000002da : MUXCY
    port map (
      CI => blk00000003_sig000003bf,
      DI => blk00000003_sig000003bc,
      S => blk00000003_sig000003c0,
      O => blk00000003_sig000003d1
    );
  blk00000003_blk000002d9 : MUXCY
    port map (
      CI => blk00000003_sig000003ce,
      DI => blk00000003_sig000003b7,
      S => blk00000003_sig000003cf,
      O => blk00000003_sig000003cb
    );
  blk00000003_blk000002d8 : MUXCY
    port map (
      CI => blk00000003_sig000003cb,
      DI => blk00000003_sig000003b8,
      S => blk00000003_sig000003cc,
      O => blk00000003_sig000003c8
    );
  blk00000003_blk000002d7 : MUXCY
    port map (
      CI => blk00000003_sig000003c8,
      DI => blk00000003_sig000003b9,
      S => blk00000003_sig000003c9,
      O => blk00000003_sig000003c5
    );
  blk00000003_blk000002d6 : MUXCY
    port map (
      CI => blk00000003_sig000003c5,
      DI => blk00000003_sig000003ba,
      S => blk00000003_sig000003c6,
      O => blk00000003_sig000003c2
    );
  blk00000003_blk000002d5 : MUXCY
    port map (
      CI => blk00000003_sig000003c2,
      DI => blk00000003_sig000003bb,
      S => blk00000003_sig000003c3,
      O => blk00000003_sig000003bf
    );
  blk00000003_blk000002d4 : XORCY
    port map (
      CI => blk00000003_sig000003ce,
      LI => blk00000003_sig000003cf,
      O => blk00000003_sig000003d0
    );
  blk00000003_blk000002d3 : XORCY
    port map (
      CI => blk00000003_sig000003cb,
      LI => blk00000003_sig000003cc,
      O => blk00000003_sig000003cd
    );
  blk00000003_blk000002d2 : XORCY
    port map (
      CI => blk00000003_sig000003c8,
      LI => blk00000003_sig000003c9,
      O => blk00000003_sig000003ca
    );
  blk00000003_blk000002d1 : XORCY
    port map (
      CI => blk00000003_sig000003c5,
      LI => blk00000003_sig000003c6,
      O => blk00000003_sig000003c7
    );
  blk00000003_blk000002d0 : XORCY
    port map (
      CI => blk00000003_sig000003c2,
      LI => blk00000003_sig000003c3,
      O => blk00000003_sig000003c4
    );
  blk00000003_blk000002cf : XORCY
    port map (
      CI => blk00000003_sig000003bf,
      LI => blk00000003_sig000003c0,
      O => blk00000003_sig000003c1
    );
  blk00000003_blk000002ce : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003b2,
      Q => blk00000003_sig000003be
    );
  blk00000003_blk000002cd : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003a2,
      Q => blk00000003_sig000003bd
    );
  blk00000003_blk000002cc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003a5,
      Q => blk00000003_sig000003bc
    );
  blk00000003_blk000002cb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003a8,
      Q => blk00000003_sig000003bb
    );
  blk00000003_blk000002ca : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003ab,
      Q => blk00000003_sig000003ba
    );
  blk00000003_blk000002c9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003ae,
      Q => blk00000003_sig000003b9
    );
  blk00000003_blk000002c8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003b1,
      Q => blk00000003_sig000003b8
    );
  blk00000003_blk000002c7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000003b5,
      Q => blk00000003_sig000003b7
    );
  blk00000003_blk000002c6 : MUXCY
    port map (
      CI => blk00000003_sig000003b3,
      DI => blk00000003_sig000003b6,
      S => blk00000003_sig000003b4,
      O => blk00000003_sig000003af
    );
  blk00000003_blk000002c5 : XORCY
    port map (
      CI => blk00000003_sig000003b3,
      LI => blk00000003_sig000003b4,
      O => blk00000003_sig000003b5
    );
  blk00000003_blk000002c4 : MUXCY
    port map (
      CI => blk00000003_sig000003a0,
      DI => blk00000003_sig0000039d,
      S => blk00000003_sig000003a1,
      O => blk00000003_sig000003b2
    );
  blk00000003_blk000002c3 : MUXCY
    port map (
      CI => blk00000003_sig000003af,
      DI => blk00000003_sig00000398,
      S => blk00000003_sig000003b0,
      O => blk00000003_sig000003ac
    );
  blk00000003_blk000002c2 : MUXCY
    port map (
      CI => blk00000003_sig000003ac,
      DI => blk00000003_sig00000399,
      S => blk00000003_sig000003ad,
      O => blk00000003_sig000003a9
    );
  blk00000003_blk000002c1 : MUXCY
    port map (
      CI => blk00000003_sig000003a9,
      DI => blk00000003_sig0000039a,
      S => blk00000003_sig000003aa,
      O => blk00000003_sig000003a6
    );
  blk00000003_blk000002c0 : MUXCY
    port map (
      CI => blk00000003_sig000003a6,
      DI => blk00000003_sig0000039b,
      S => blk00000003_sig000003a7,
      O => blk00000003_sig000003a3
    );
  blk00000003_blk000002bf : MUXCY
    port map (
      CI => blk00000003_sig000003a3,
      DI => blk00000003_sig0000039c,
      S => blk00000003_sig000003a4,
      O => blk00000003_sig000003a0
    );
  blk00000003_blk000002be : XORCY
    port map (
      CI => blk00000003_sig000003af,
      LI => blk00000003_sig000003b0,
      O => blk00000003_sig000003b1
    );
  blk00000003_blk000002bd : XORCY
    port map (
      CI => blk00000003_sig000003ac,
      LI => blk00000003_sig000003ad,
      O => blk00000003_sig000003ae
    );
  blk00000003_blk000002bc : XORCY
    port map (
      CI => blk00000003_sig000003a9,
      LI => blk00000003_sig000003aa,
      O => blk00000003_sig000003ab
    );
  blk00000003_blk000002bb : XORCY
    port map (
      CI => blk00000003_sig000003a6,
      LI => blk00000003_sig000003a7,
      O => blk00000003_sig000003a8
    );
  blk00000003_blk000002ba : XORCY
    port map (
      CI => blk00000003_sig000003a3,
      LI => blk00000003_sig000003a4,
      O => blk00000003_sig000003a5
    );
  blk00000003_blk000002b9 : XORCY
    port map (
      CI => blk00000003_sig000003a0,
      LI => blk00000003_sig000003a1,
      O => blk00000003_sig000003a2
    );
  blk00000003_blk000002b8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000393,
      Q => blk00000003_sig0000039f
    );
  blk00000003_blk000002b7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000383,
      Q => blk00000003_sig0000039e
    );
  blk00000003_blk000002b6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000386,
      Q => blk00000003_sig0000039d
    );
  blk00000003_blk000002b5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000389,
      Q => blk00000003_sig0000039c
    );
  blk00000003_blk000002b4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000038c,
      Q => blk00000003_sig0000039b
    );
  blk00000003_blk000002b3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000038f,
      Q => blk00000003_sig0000039a
    );
  blk00000003_blk000002b2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000392,
      Q => blk00000003_sig00000399
    );
  blk00000003_blk000002b1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000396,
      Q => blk00000003_sig00000398
    );
  blk00000003_blk000002b0 : MUXCY
    port map (
      CI => blk00000003_sig00000394,
      DI => blk00000003_sig00000397,
      S => blk00000003_sig00000395,
      O => blk00000003_sig00000390
    );
  blk00000003_blk000002af : XORCY
    port map (
      CI => blk00000003_sig00000394,
      LI => blk00000003_sig00000395,
      O => blk00000003_sig00000396
    );
  blk00000003_blk000002ae : MUXCY
    port map (
      CI => blk00000003_sig00000381,
      DI => blk00000003_sig0000037e,
      S => blk00000003_sig00000382,
      O => blk00000003_sig00000393
    );
  blk00000003_blk000002ad : MUXCY
    port map (
      CI => blk00000003_sig00000390,
      DI => blk00000003_sig00000379,
      S => blk00000003_sig00000391,
      O => blk00000003_sig0000038d
    );
  blk00000003_blk000002ac : MUXCY
    port map (
      CI => blk00000003_sig0000038d,
      DI => blk00000003_sig0000037a,
      S => blk00000003_sig0000038e,
      O => blk00000003_sig0000038a
    );
  blk00000003_blk000002ab : MUXCY
    port map (
      CI => blk00000003_sig0000038a,
      DI => blk00000003_sig0000037b,
      S => blk00000003_sig0000038b,
      O => blk00000003_sig00000387
    );
  blk00000003_blk000002aa : MUXCY
    port map (
      CI => blk00000003_sig00000387,
      DI => blk00000003_sig0000037c,
      S => blk00000003_sig00000388,
      O => blk00000003_sig00000384
    );
  blk00000003_blk000002a9 : MUXCY
    port map (
      CI => blk00000003_sig00000384,
      DI => blk00000003_sig0000037d,
      S => blk00000003_sig00000385,
      O => blk00000003_sig00000381
    );
  blk00000003_blk000002a8 : XORCY
    port map (
      CI => blk00000003_sig00000390,
      LI => blk00000003_sig00000391,
      O => blk00000003_sig00000392
    );
  blk00000003_blk000002a7 : XORCY
    port map (
      CI => blk00000003_sig0000038d,
      LI => blk00000003_sig0000038e,
      O => blk00000003_sig0000038f
    );
  blk00000003_blk000002a6 : XORCY
    port map (
      CI => blk00000003_sig0000038a,
      LI => blk00000003_sig0000038b,
      O => blk00000003_sig0000038c
    );
  blk00000003_blk000002a5 : XORCY
    port map (
      CI => blk00000003_sig00000387,
      LI => blk00000003_sig00000388,
      O => blk00000003_sig00000389
    );
  blk00000003_blk000002a4 : XORCY
    port map (
      CI => blk00000003_sig00000384,
      LI => blk00000003_sig00000385,
      O => blk00000003_sig00000386
    );
  blk00000003_blk000002a3 : XORCY
    port map (
      CI => blk00000003_sig00000381,
      LI => blk00000003_sig00000382,
      O => blk00000003_sig00000383
    );
  blk00000003_blk000002a2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000374,
      Q => blk00000003_sig00000380
    );
  blk00000003_blk000002a1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000364,
      Q => blk00000003_sig0000037f
    );
  blk00000003_blk000002a0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000367,
      Q => blk00000003_sig0000037e
    );
  blk00000003_blk0000029f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000036a,
      Q => blk00000003_sig0000037d
    );
  blk00000003_blk0000029e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000036d,
      Q => blk00000003_sig0000037c
    );
  blk00000003_blk0000029d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000370,
      Q => blk00000003_sig0000037b
    );
  blk00000003_blk0000029c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000373,
      Q => blk00000003_sig0000037a
    );
  blk00000003_blk0000029b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000377,
      Q => blk00000003_sig00000379
    );
  blk00000003_blk0000029a : MUXCY
    port map (
      CI => blk00000003_sig00000375,
      DI => blk00000003_sig00000378,
      S => blk00000003_sig00000376,
      O => blk00000003_sig00000371
    );
  blk00000003_blk00000299 : XORCY
    port map (
      CI => blk00000003_sig00000375,
      LI => blk00000003_sig00000376,
      O => blk00000003_sig00000377
    );
  blk00000003_blk00000298 : MUXCY
    port map (
      CI => blk00000003_sig00000362,
      DI => blk00000003_sig0000035f,
      S => blk00000003_sig00000363,
      O => blk00000003_sig00000374
    );
  blk00000003_blk00000297 : MUXCY
    port map (
      CI => blk00000003_sig00000371,
      DI => blk00000003_sig0000035a,
      S => blk00000003_sig00000372,
      O => blk00000003_sig0000036e
    );
  blk00000003_blk00000296 : MUXCY
    port map (
      CI => blk00000003_sig0000036e,
      DI => blk00000003_sig0000035b,
      S => blk00000003_sig0000036f,
      O => blk00000003_sig0000036b
    );
  blk00000003_blk00000295 : MUXCY
    port map (
      CI => blk00000003_sig0000036b,
      DI => blk00000003_sig0000035c,
      S => blk00000003_sig0000036c,
      O => blk00000003_sig00000368
    );
  blk00000003_blk00000294 : MUXCY
    port map (
      CI => blk00000003_sig00000368,
      DI => blk00000003_sig0000035d,
      S => blk00000003_sig00000369,
      O => blk00000003_sig00000365
    );
  blk00000003_blk00000293 : MUXCY
    port map (
      CI => blk00000003_sig00000365,
      DI => blk00000003_sig0000035e,
      S => blk00000003_sig00000366,
      O => blk00000003_sig00000362
    );
  blk00000003_blk00000292 : XORCY
    port map (
      CI => blk00000003_sig00000371,
      LI => blk00000003_sig00000372,
      O => blk00000003_sig00000373
    );
  blk00000003_blk00000291 : XORCY
    port map (
      CI => blk00000003_sig0000036e,
      LI => blk00000003_sig0000036f,
      O => blk00000003_sig00000370
    );
  blk00000003_blk00000290 : XORCY
    port map (
      CI => blk00000003_sig0000036b,
      LI => blk00000003_sig0000036c,
      O => blk00000003_sig0000036d
    );
  blk00000003_blk0000028f : XORCY
    port map (
      CI => blk00000003_sig00000368,
      LI => blk00000003_sig00000369,
      O => blk00000003_sig0000036a
    );
  blk00000003_blk0000028e : XORCY
    port map (
      CI => blk00000003_sig00000365,
      LI => blk00000003_sig00000366,
      O => blk00000003_sig00000367
    );
  blk00000003_blk0000028d : XORCY
    port map (
      CI => blk00000003_sig00000362,
      LI => blk00000003_sig00000363,
      O => blk00000003_sig00000364
    );
  blk00000003_blk0000028c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000355,
      Q => blk00000003_sig00000361
    );
  blk00000003_blk0000028b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000345,
      Q => blk00000003_sig00000360
    );
  blk00000003_blk0000028a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000348,
      Q => blk00000003_sig0000035f
    );
  blk00000003_blk00000289 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000034b,
      Q => blk00000003_sig0000035e
    );
  blk00000003_blk00000288 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000034e,
      Q => blk00000003_sig0000035d
    );
  blk00000003_blk00000287 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000351,
      Q => blk00000003_sig0000035c
    );
  blk00000003_blk00000286 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000354,
      Q => blk00000003_sig0000035b
    );
  blk00000003_blk00000285 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000358,
      Q => blk00000003_sig0000035a
    );
  blk00000003_blk00000284 : MUXCY
    port map (
      CI => blk00000003_sig00000356,
      DI => blk00000003_sig00000359,
      S => blk00000003_sig00000357,
      O => blk00000003_sig00000352
    );
  blk00000003_blk00000283 : XORCY
    port map (
      CI => blk00000003_sig00000356,
      LI => blk00000003_sig00000357,
      O => blk00000003_sig00000358
    );
  blk00000003_blk00000282 : MUXCY
    port map (
      CI => blk00000003_sig00000343,
      DI => blk00000003_sig00000340,
      S => blk00000003_sig00000344,
      O => blk00000003_sig00000355
    );
  blk00000003_blk00000281 : MUXCY
    port map (
      CI => blk00000003_sig00000352,
      DI => blk00000003_sig0000033b,
      S => blk00000003_sig00000353,
      O => blk00000003_sig0000034f
    );
  blk00000003_blk00000280 : MUXCY
    port map (
      CI => blk00000003_sig0000034f,
      DI => blk00000003_sig0000033c,
      S => blk00000003_sig00000350,
      O => blk00000003_sig0000034c
    );
  blk00000003_blk0000027f : MUXCY
    port map (
      CI => blk00000003_sig0000034c,
      DI => blk00000003_sig0000033d,
      S => blk00000003_sig0000034d,
      O => blk00000003_sig00000349
    );
  blk00000003_blk0000027e : MUXCY
    port map (
      CI => blk00000003_sig00000349,
      DI => blk00000003_sig0000033e,
      S => blk00000003_sig0000034a,
      O => blk00000003_sig00000346
    );
  blk00000003_blk0000027d : MUXCY
    port map (
      CI => blk00000003_sig00000346,
      DI => blk00000003_sig0000033f,
      S => blk00000003_sig00000347,
      O => blk00000003_sig00000343
    );
  blk00000003_blk0000027c : XORCY
    port map (
      CI => blk00000003_sig00000352,
      LI => blk00000003_sig00000353,
      O => blk00000003_sig00000354
    );
  blk00000003_blk0000027b : XORCY
    port map (
      CI => blk00000003_sig0000034f,
      LI => blk00000003_sig00000350,
      O => blk00000003_sig00000351
    );
  blk00000003_blk0000027a : XORCY
    port map (
      CI => blk00000003_sig0000034c,
      LI => blk00000003_sig0000034d,
      O => blk00000003_sig0000034e
    );
  blk00000003_blk00000279 : XORCY
    port map (
      CI => blk00000003_sig00000349,
      LI => blk00000003_sig0000034a,
      O => blk00000003_sig0000034b
    );
  blk00000003_blk00000278 : XORCY
    port map (
      CI => blk00000003_sig00000346,
      LI => blk00000003_sig00000347,
      O => blk00000003_sig00000348
    );
  blk00000003_blk00000277 : XORCY
    port map (
      CI => blk00000003_sig00000343,
      LI => blk00000003_sig00000344,
      O => blk00000003_sig00000345
    );
  blk00000003_blk00000276 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000336,
      Q => blk00000003_sig00000342
    );
  blk00000003_blk00000275 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000326,
      Q => blk00000003_sig00000341
    );
  blk00000003_blk00000274 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000329,
      Q => blk00000003_sig00000340
    );
  blk00000003_blk00000273 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000032c,
      Q => blk00000003_sig0000033f
    );
  blk00000003_blk00000272 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000032f,
      Q => blk00000003_sig0000033e
    );
  blk00000003_blk00000271 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000332,
      Q => blk00000003_sig0000033d
    );
  blk00000003_blk00000270 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000335,
      Q => blk00000003_sig0000033c
    );
  blk00000003_blk0000026f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000339,
      Q => blk00000003_sig0000033b
    );
  blk00000003_blk0000026e : MUXCY
    port map (
      CI => blk00000003_sig00000337,
      DI => blk00000003_sig0000033a,
      S => blk00000003_sig00000338,
      O => blk00000003_sig00000333
    );
  blk00000003_blk0000026d : XORCY
    port map (
      CI => blk00000003_sig00000337,
      LI => blk00000003_sig00000338,
      O => blk00000003_sig00000339
    );
  blk00000003_blk0000026c : MUXCY
    port map (
      CI => blk00000003_sig00000324,
      DI => blk00000003_sig00000321,
      S => blk00000003_sig00000325,
      O => blk00000003_sig00000336
    );
  blk00000003_blk0000026b : MUXCY
    port map (
      CI => blk00000003_sig00000333,
      DI => blk00000003_sig0000031c,
      S => blk00000003_sig00000334,
      O => blk00000003_sig00000330
    );
  blk00000003_blk0000026a : MUXCY
    port map (
      CI => blk00000003_sig00000330,
      DI => blk00000003_sig0000031d,
      S => blk00000003_sig00000331,
      O => blk00000003_sig0000032d
    );
  blk00000003_blk00000269 : MUXCY
    port map (
      CI => blk00000003_sig0000032d,
      DI => blk00000003_sig0000031e,
      S => blk00000003_sig0000032e,
      O => blk00000003_sig0000032a
    );
  blk00000003_blk00000268 : MUXCY
    port map (
      CI => blk00000003_sig0000032a,
      DI => blk00000003_sig0000031f,
      S => blk00000003_sig0000032b,
      O => blk00000003_sig00000327
    );
  blk00000003_blk00000267 : MUXCY
    port map (
      CI => blk00000003_sig00000327,
      DI => blk00000003_sig00000320,
      S => blk00000003_sig00000328,
      O => blk00000003_sig00000324
    );
  blk00000003_blk00000266 : XORCY
    port map (
      CI => blk00000003_sig00000333,
      LI => blk00000003_sig00000334,
      O => blk00000003_sig00000335
    );
  blk00000003_blk00000265 : XORCY
    port map (
      CI => blk00000003_sig00000330,
      LI => blk00000003_sig00000331,
      O => blk00000003_sig00000332
    );
  blk00000003_blk00000264 : XORCY
    port map (
      CI => blk00000003_sig0000032d,
      LI => blk00000003_sig0000032e,
      O => blk00000003_sig0000032f
    );
  blk00000003_blk00000263 : XORCY
    port map (
      CI => blk00000003_sig0000032a,
      LI => blk00000003_sig0000032b,
      O => blk00000003_sig0000032c
    );
  blk00000003_blk00000262 : XORCY
    port map (
      CI => blk00000003_sig00000327,
      LI => blk00000003_sig00000328,
      O => blk00000003_sig00000329
    );
  blk00000003_blk00000261 : XORCY
    port map (
      CI => blk00000003_sig00000324,
      LI => blk00000003_sig00000325,
      O => blk00000003_sig00000326
    );
  blk00000003_blk00000260 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000317,
      Q => blk00000003_sig00000323
    );
  blk00000003_blk0000025f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000307,
      Q => blk00000003_sig00000322
    );
  blk00000003_blk0000025e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000030a,
      Q => blk00000003_sig00000321
    );
  blk00000003_blk0000025d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000030d,
      Q => blk00000003_sig00000320
    );
  blk00000003_blk0000025c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000310,
      Q => blk00000003_sig0000031f
    );
  blk00000003_blk0000025b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000313,
      Q => blk00000003_sig0000031e
    );
  blk00000003_blk0000025a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000316,
      Q => blk00000003_sig0000031d
    );
  blk00000003_blk00000259 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000031a,
      Q => blk00000003_sig0000031c
    );
  blk00000003_blk00000258 : MUXCY
    port map (
      CI => blk00000003_sig00000318,
      DI => blk00000003_sig0000031b,
      S => blk00000003_sig00000319,
      O => blk00000003_sig00000314
    );
  blk00000003_blk00000257 : XORCY
    port map (
      CI => blk00000003_sig00000318,
      LI => blk00000003_sig00000319,
      O => blk00000003_sig0000031a
    );
  blk00000003_blk00000256 : MUXCY
    port map (
      CI => blk00000003_sig00000305,
      DI => blk00000003_sig00000302,
      S => blk00000003_sig00000306,
      O => blk00000003_sig00000317
    );
  blk00000003_blk00000255 : MUXCY
    port map (
      CI => blk00000003_sig00000314,
      DI => blk00000003_sig000002fd,
      S => blk00000003_sig00000315,
      O => blk00000003_sig00000311
    );
  blk00000003_blk00000254 : MUXCY
    port map (
      CI => blk00000003_sig00000311,
      DI => blk00000003_sig000002fe,
      S => blk00000003_sig00000312,
      O => blk00000003_sig0000030e
    );
  blk00000003_blk00000253 : MUXCY
    port map (
      CI => blk00000003_sig0000030e,
      DI => blk00000003_sig000002ff,
      S => blk00000003_sig0000030f,
      O => blk00000003_sig0000030b
    );
  blk00000003_blk00000252 : MUXCY
    port map (
      CI => blk00000003_sig0000030b,
      DI => blk00000003_sig00000300,
      S => blk00000003_sig0000030c,
      O => blk00000003_sig00000308
    );
  blk00000003_blk00000251 : MUXCY
    port map (
      CI => blk00000003_sig00000308,
      DI => blk00000003_sig00000301,
      S => blk00000003_sig00000309,
      O => blk00000003_sig00000305
    );
  blk00000003_blk00000250 : XORCY
    port map (
      CI => blk00000003_sig00000314,
      LI => blk00000003_sig00000315,
      O => blk00000003_sig00000316
    );
  blk00000003_blk0000024f : XORCY
    port map (
      CI => blk00000003_sig00000311,
      LI => blk00000003_sig00000312,
      O => blk00000003_sig00000313
    );
  blk00000003_blk0000024e : XORCY
    port map (
      CI => blk00000003_sig0000030e,
      LI => blk00000003_sig0000030f,
      O => blk00000003_sig00000310
    );
  blk00000003_blk0000024d : XORCY
    port map (
      CI => blk00000003_sig0000030b,
      LI => blk00000003_sig0000030c,
      O => blk00000003_sig0000030d
    );
  blk00000003_blk0000024c : XORCY
    port map (
      CI => blk00000003_sig00000308,
      LI => blk00000003_sig00000309,
      O => blk00000003_sig0000030a
    );
  blk00000003_blk0000024b : XORCY
    port map (
      CI => blk00000003_sig00000305,
      LI => blk00000003_sig00000306,
      O => blk00000003_sig00000307
    );
  blk00000003_blk0000024a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002f8,
      Q => blk00000003_sig00000304
    );
  blk00000003_blk00000249 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002e8,
      Q => blk00000003_sig00000303
    );
  blk00000003_blk00000248 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002eb,
      Q => blk00000003_sig00000302
    );
  blk00000003_blk00000247 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002ee,
      Q => blk00000003_sig00000301
    );
  blk00000003_blk00000246 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002f1,
      Q => blk00000003_sig00000300
    );
  blk00000003_blk00000245 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002f4,
      Q => blk00000003_sig000002ff
    );
  blk00000003_blk00000244 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002f7,
      Q => blk00000003_sig000002fe
    );
  blk00000003_blk00000243 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002fb,
      Q => blk00000003_sig000002fd
    );
  blk00000003_blk00000242 : MUXCY
    port map (
      CI => blk00000003_sig000002f9,
      DI => blk00000003_sig000002fc,
      S => blk00000003_sig000002fa,
      O => blk00000003_sig000002f5
    );
  blk00000003_blk00000241 : XORCY
    port map (
      CI => blk00000003_sig000002f9,
      LI => blk00000003_sig000002fa,
      O => blk00000003_sig000002fb
    );
  blk00000003_blk00000240 : MUXCY
    port map (
      CI => blk00000003_sig000002e6,
      DI => blk00000003_sig000002e3,
      S => blk00000003_sig000002e7,
      O => blk00000003_sig000002f8
    );
  blk00000003_blk0000023f : MUXCY
    port map (
      CI => blk00000003_sig000002f5,
      DI => blk00000003_sig000002de,
      S => blk00000003_sig000002f6,
      O => blk00000003_sig000002f2
    );
  blk00000003_blk0000023e : MUXCY
    port map (
      CI => blk00000003_sig000002f2,
      DI => blk00000003_sig000002df,
      S => blk00000003_sig000002f3,
      O => blk00000003_sig000002ef
    );
  blk00000003_blk0000023d : MUXCY
    port map (
      CI => blk00000003_sig000002ef,
      DI => blk00000003_sig000002e0,
      S => blk00000003_sig000002f0,
      O => blk00000003_sig000002ec
    );
  blk00000003_blk0000023c : MUXCY
    port map (
      CI => blk00000003_sig000002ec,
      DI => blk00000003_sig000002e1,
      S => blk00000003_sig000002ed,
      O => blk00000003_sig000002e9
    );
  blk00000003_blk0000023b : MUXCY
    port map (
      CI => blk00000003_sig000002e9,
      DI => blk00000003_sig000002e2,
      S => blk00000003_sig000002ea,
      O => blk00000003_sig000002e6
    );
  blk00000003_blk0000023a : XORCY
    port map (
      CI => blk00000003_sig000002f5,
      LI => blk00000003_sig000002f6,
      O => blk00000003_sig000002f7
    );
  blk00000003_blk00000239 : XORCY
    port map (
      CI => blk00000003_sig000002f2,
      LI => blk00000003_sig000002f3,
      O => blk00000003_sig000002f4
    );
  blk00000003_blk00000238 : XORCY
    port map (
      CI => blk00000003_sig000002ef,
      LI => blk00000003_sig000002f0,
      O => blk00000003_sig000002f1
    );
  blk00000003_blk00000237 : XORCY
    port map (
      CI => blk00000003_sig000002ec,
      LI => blk00000003_sig000002ed,
      O => blk00000003_sig000002ee
    );
  blk00000003_blk00000236 : XORCY
    port map (
      CI => blk00000003_sig000002e9,
      LI => blk00000003_sig000002ea,
      O => blk00000003_sig000002eb
    );
  blk00000003_blk00000235 : XORCY
    port map (
      CI => blk00000003_sig000002e6,
      LI => blk00000003_sig000002e7,
      O => blk00000003_sig000002e8
    );
  blk00000003_blk00000234 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002d9,
      Q => blk00000003_sig000002e5
    );
  blk00000003_blk00000233 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002c9,
      Q => blk00000003_sig000002e4
    );
  blk00000003_blk00000232 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002cc,
      Q => blk00000003_sig000002e3
    );
  blk00000003_blk00000231 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002cf,
      Q => blk00000003_sig000002e2
    );
  blk00000003_blk00000230 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002d2,
      Q => blk00000003_sig000002e1
    );
  blk00000003_blk0000022f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002d5,
      Q => blk00000003_sig000002e0
    );
  blk00000003_blk0000022e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002d8,
      Q => blk00000003_sig000002df
    );
  blk00000003_blk0000022d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002dc,
      Q => blk00000003_sig000002de
    );
  blk00000003_blk0000022c : MUXCY
    port map (
      CI => blk00000003_sig000002da,
      DI => blk00000003_sig000002dd,
      S => blk00000003_sig000002db,
      O => blk00000003_sig000002d6
    );
  blk00000003_blk0000022b : XORCY
    port map (
      CI => blk00000003_sig000002da,
      LI => blk00000003_sig000002db,
      O => blk00000003_sig000002dc
    );
  blk00000003_blk0000022a : MUXCY
    port map (
      CI => blk00000003_sig000002c7,
      DI => blk00000003_sig000002c4,
      S => blk00000003_sig000002c8,
      O => blk00000003_sig000002d9
    );
  blk00000003_blk00000229 : MUXCY
    port map (
      CI => blk00000003_sig000002d6,
      DI => blk00000003_sig000002bf,
      S => blk00000003_sig000002d7,
      O => blk00000003_sig000002d3
    );
  blk00000003_blk00000228 : MUXCY
    port map (
      CI => blk00000003_sig000002d3,
      DI => blk00000003_sig000002c0,
      S => blk00000003_sig000002d4,
      O => blk00000003_sig000002d0
    );
  blk00000003_blk00000227 : MUXCY
    port map (
      CI => blk00000003_sig000002d0,
      DI => blk00000003_sig000002c1,
      S => blk00000003_sig000002d1,
      O => blk00000003_sig000002cd
    );
  blk00000003_blk00000226 : MUXCY
    port map (
      CI => blk00000003_sig000002cd,
      DI => blk00000003_sig000002c2,
      S => blk00000003_sig000002ce,
      O => blk00000003_sig000002ca
    );
  blk00000003_blk00000225 : MUXCY
    port map (
      CI => blk00000003_sig000002ca,
      DI => blk00000003_sig000002c3,
      S => blk00000003_sig000002cb,
      O => blk00000003_sig000002c7
    );
  blk00000003_blk00000224 : XORCY
    port map (
      CI => blk00000003_sig000002d6,
      LI => blk00000003_sig000002d7,
      O => blk00000003_sig000002d8
    );
  blk00000003_blk00000223 : XORCY
    port map (
      CI => blk00000003_sig000002d3,
      LI => blk00000003_sig000002d4,
      O => blk00000003_sig000002d5
    );
  blk00000003_blk00000222 : XORCY
    port map (
      CI => blk00000003_sig000002d0,
      LI => blk00000003_sig000002d1,
      O => blk00000003_sig000002d2
    );
  blk00000003_blk00000221 : XORCY
    port map (
      CI => blk00000003_sig000002cd,
      LI => blk00000003_sig000002ce,
      O => blk00000003_sig000002cf
    );
  blk00000003_blk00000220 : XORCY
    port map (
      CI => blk00000003_sig000002ca,
      LI => blk00000003_sig000002cb,
      O => blk00000003_sig000002cc
    );
  blk00000003_blk0000021f : XORCY
    port map (
      CI => blk00000003_sig000002c7,
      LI => blk00000003_sig000002c8,
      O => blk00000003_sig000002c9
    );
  blk00000003_blk0000021e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002ba,
      Q => blk00000003_sig000002c6
    );
  blk00000003_blk0000021d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002aa,
      Q => blk00000003_sig000002c5
    );
  blk00000003_blk0000021c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002ad,
      Q => blk00000003_sig000002c4
    );
  blk00000003_blk0000021b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002b0,
      Q => blk00000003_sig000002c3
    );
  blk00000003_blk0000021a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002b3,
      Q => blk00000003_sig000002c2
    );
  blk00000003_blk00000219 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002b6,
      Q => blk00000003_sig000002c1
    );
  blk00000003_blk00000218 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002b9,
      Q => blk00000003_sig000002c0
    );
  blk00000003_blk00000217 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000002bd,
      Q => blk00000003_sig000002bf
    );
  blk00000003_blk00000216 : MUXCY
    port map (
      CI => blk00000003_sig000002bb,
      DI => blk00000003_sig000002be,
      S => blk00000003_sig000002bc,
      O => blk00000003_sig000002b7
    );
  blk00000003_blk00000215 : XORCY
    port map (
      CI => blk00000003_sig000002bb,
      LI => blk00000003_sig000002bc,
      O => blk00000003_sig000002bd
    );
  blk00000003_blk00000214 : MUXCY
    port map (
      CI => blk00000003_sig000002a8,
      DI => blk00000003_sig000002a5,
      S => blk00000003_sig000002a9,
      O => blk00000003_sig000002ba
    );
  blk00000003_blk00000213 : MUXCY
    port map (
      CI => blk00000003_sig000002b7,
      DI => blk00000003_sig000002a0,
      S => blk00000003_sig000002b8,
      O => blk00000003_sig000002b4
    );
  blk00000003_blk00000212 : MUXCY
    port map (
      CI => blk00000003_sig000002b4,
      DI => blk00000003_sig000002a1,
      S => blk00000003_sig000002b5,
      O => blk00000003_sig000002b1
    );
  blk00000003_blk00000211 : MUXCY
    port map (
      CI => blk00000003_sig000002b1,
      DI => blk00000003_sig000002a2,
      S => blk00000003_sig000002b2,
      O => blk00000003_sig000002ae
    );
  blk00000003_blk00000210 : MUXCY
    port map (
      CI => blk00000003_sig000002ae,
      DI => blk00000003_sig000002a3,
      S => blk00000003_sig000002af,
      O => blk00000003_sig000002ab
    );
  blk00000003_blk0000020f : MUXCY
    port map (
      CI => blk00000003_sig000002ab,
      DI => blk00000003_sig000002a4,
      S => blk00000003_sig000002ac,
      O => blk00000003_sig000002a8
    );
  blk00000003_blk0000020e : XORCY
    port map (
      CI => blk00000003_sig000002b7,
      LI => blk00000003_sig000002b8,
      O => blk00000003_sig000002b9
    );
  blk00000003_blk0000020d : XORCY
    port map (
      CI => blk00000003_sig000002b4,
      LI => blk00000003_sig000002b5,
      O => blk00000003_sig000002b6
    );
  blk00000003_blk0000020c : XORCY
    port map (
      CI => blk00000003_sig000002b1,
      LI => blk00000003_sig000002b2,
      O => blk00000003_sig000002b3
    );
  blk00000003_blk0000020b : XORCY
    port map (
      CI => blk00000003_sig000002ae,
      LI => blk00000003_sig000002af,
      O => blk00000003_sig000002b0
    );
  blk00000003_blk0000020a : XORCY
    port map (
      CI => blk00000003_sig000002ab,
      LI => blk00000003_sig000002ac,
      O => blk00000003_sig000002ad
    );
  blk00000003_blk00000209 : XORCY
    port map (
      CI => blk00000003_sig000002a8,
      LI => blk00000003_sig000002a9,
      O => blk00000003_sig000002aa
    );
  blk00000003_blk00000208 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000029b,
      Q => blk00000003_sig000002a7
    );
  blk00000003_blk00000207 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000028b,
      Q => blk00000003_sig000002a6
    );
  blk00000003_blk00000206 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000028e,
      Q => blk00000003_sig000002a5
    );
  blk00000003_blk00000205 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000291,
      Q => blk00000003_sig000002a4
    );
  blk00000003_blk00000204 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000294,
      Q => blk00000003_sig000002a3
    );
  blk00000003_blk00000203 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000297,
      Q => blk00000003_sig000002a2
    );
  blk00000003_blk00000202 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000029a,
      Q => blk00000003_sig000002a1
    );
  blk00000003_blk00000201 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000029e,
      Q => blk00000003_sig000002a0
    );
  blk00000003_blk00000200 : MUXCY
    port map (
      CI => blk00000003_sig0000029c,
      DI => blk00000003_sig0000029f,
      S => blk00000003_sig0000029d,
      O => blk00000003_sig00000298
    );
  blk00000003_blk000001ff : XORCY
    port map (
      CI => blk00000003_sig0000029c,
      LI => blk00000003_sig0000029d,
      O => blk00000003_sig0000029e
    );
  blk00000003_blk000001fe : MUXCY
    port map (
      CI => blk00000003_sig00000289,
      DI => blk00000003_sig00000286,
      S => blk00000003_sig0000028a,
      O => blk00000003_sig0000029b
    );
  blk00000003_blk000001fd : MUXCY
    port map (
      CI => blk00000003_sig00000298,
      DI => blk00000003_sig00000281,
      S => blk00000003_sig00000299,
      O => blk00000003_sig00000295
    );
  blk00000003_blk000001fc : MUXCY
    port map (
      CI => blk00000003_sig00000295,
      DI => blk00000003_sig00000282,
      S => blk00000003_sig00000296,
      O => blk00000003_sig00000292
    );
  blk00000003_blk000001fb : MUXCY
    port map (
      CI => blk00000003_sig00000292,
      DI => blk00000003_sig00000283,
      S => blk00000003_sig00000293,
      O => blk00000003_sig0000028f
    );
  blk00000003_blk000001fa : MUXCY
    port map (
      CI => blk00000003_sig0000028f,
      DI => blk00000003_sig00000284,
      S => blk00000003_sig00000290,
      O => blk00000003_sig0000028c
    );
  blk00000003_blk000001f9 : MUXCY
    port map (
      CI => blk00000003_sig0000028c,
      DI => blk00000003_sig00000285,
      S => blk00000003_sig0000028d,
      O => blk00000003_sig00000289
    );
  blk00000003_blk000001f8 : XORCY
    port map (
      CI => blk00000003_sig00000298,
      LI => blk00000003_sig00000299,
      O => blk00000003_sig0000029a
    );
  blk00000003_blk000001f7 : XORCY
    port map (
      CI => blk00000003_sig00000295,
      LI => blk00000003_sig00000296,
      O => blk00000003_sig00000297
    );
  blk00000003_blk000001f6 : XORCY
    port map (
      CI => blk00000003_sig00000292,
      LI => blk00000003_sig00000293,
      O => blk00000003_sig00000294
    );
  blk00000003_blk000001f5 : XORCY
    port map (
      CI => blk00000003_sig0000028f,
      LI => blk00000003_sig00000290,
      O => blk00000003_sig00000291
    );
  blk00000003_blk000001f4 : XORCY
    port map (
      CI => blk00000003_sig0000028c,
      LI => blk00000003_sig0000028d,
      O => blk00000003_sig0000028e
    );
  blk00000003_blk000001f3 : XORCY
    port map (
      CI => blk00000003_sig00000289,
      LI => blk00000003_sig0000028a,
      O => blk00000003_sig0000028b
    );
  blk00000003_blk000001f2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000027c,
      Q => blk00000003_sig00000288
    );
  blk00000003_blk000001f1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000026c,
      Q => blk00000003_sig00000287
    );
  blk00000003_blk000001f0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000026f,
      Q => blk00000003_sig00000286
    );
  blk00000003_blk000001ef : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000272,
      Q => blk00000003_sig00000285
    );
  blk00000003_blk000001ee : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000275,
      Q => blk00000003_sig00000284
    );
  blk00000003_blk000001ed : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000278,
      Q => blk00000003_sig00000283
    );
  blk00000003_blk000001ec : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000027b,
      Q => blk00000003_sig00000282
    );
  blk00000003_blk000001eb : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000027f,
      Q => blk00000003_sig00000281
    );
  blk00000003_blk000001ea : MUXCY
    port map (
      CI => blk00000003_sig0000027d,
      DI => blk00000003_sig00000280,
      S => blk00000003_sig0000027e,
      O => blk00000003_sig00000279
    );
  blk00000003_blk000001e9 : XORCY
    port map (
      CI => blk00000003_sig0000027d,
      LI => blk00000003_sig0000027e,
      O => blk00000003_sig0000027f
    );
  blk00000003_blk000001e8 : MUXCY
    port map (
      CI => blk00000003_sig0000026a,
      DI => blk00000003_sig00000268,
      S => blk00000003_sig0000026b,
      O => blk00000003_sig0000027c
    );
  blk00000003_blk000001e7 : MUXCY
    port map (
      CI => blk00000003_sig00000279,
      DI => blk00000003_sig00000263,
      S => blk00000003_sig0000027a,
      O => blk00000003_sig00000276
    );
  blk00000003_blk000001e6 : MUXCY
    port map (
      CI => blk00000003_sig00000276,
      DI => blk00000003_sig00000264,
      S => blk00000003_sig00000277,
      O => blk00000003_sig00000273
    );
  blk00000003_blk000001e5 : MUXCY
    port map (
      CI => blk00000003_sig00000273,
      DI => blk00000003_sig00000265,
      S => blk00000003_sig00000274,
      O => blk00000003_sig00000270
    );
  blk00000003_blk000001e4 : MUXCY
    port map (
      CI => blk00000003_sig00000270,
      DI => blk00000003_sig00000266,
      S => blk00000003_sig00000271,
      O => blk00000003_sig0000026d
    );
  blk00000003_blk000001e3 : MUXCY
    port map (
      CI => blk00000003_sig0000026d,
      DI => blk00000003_sig00000267,
      S => blk00000003_sig0000026e,
      O => blk00000003_sig0000026a
    );
  blk00000003_blk000001e2 : XORCY
    port map (
      CI => blk00000003_sig00000279,
      LI => blk00000003_sig0000027a,
      O => blk00000003_sig0000027b
    );
  blk00000003_blk000001e1 : XORCY
    port map (
      CI => blk00000003_sig00000276,
      LI => blk00000003_sig00000277,
      O => blk00000003_sig00000278
    );
  blk00000003_blk000001e0 : XORCY
    port map (
      CI => blk00000003_sig00000273,
      LI => blk00000003_sig00000274,
      O => blk00000003_sig00000275
    );
  blk00000003_blk000001df : XORCY
    port map (
      CI => blk00000003_sig00000270,
      LI => blk00000003_sig00000271,
      O => blk00000003_sig00000272
    );
  blk00000003_blk000001de : XORCY
    port map (
      CI => blk00000003_sig0000026d,
      LI => blk00000003_sig0000026e,
      O => blk00000003_sig0000026f
    );
  blk00000003_blk000001dd : XORCY
    port map (
      CI => blk00000003_sig0000026a,
      LI => blk00000003_sig0000026b,
      O => blk00000003_sig0000026c
    );
  blk00000003_blk000001dc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000025e,
      Q => blk00000003_sig00000269
    );
  blk00000003_blk000001db : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000024e,
      Q => blk00000003_sig0000008e
    );
  blk00000003_blk000001da : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000251,
      Q => blk00000003_sig00000268
    );
  blk00000003_blk000001d9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000254,
      Q => blk00000003_sig00000267
    );
  blk00000003_blk000001d8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000257,
      Q => blk00000003_sig00000266
    );
  blk00000003_blk000001d7 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000025a,
      Q => blk00000003_sig00000265
    );
  blk00000003_blk000001d6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000025d,
      Q => blk00000003_sig00000264
    );
  blk00000003_blk000001d5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000261,
      Q => blk00000003_sig00000263
    );
  blk00000003_blk000001d4 : MUXCY
    port map (
      CI => blk00000003_sig0000025f,
      DI => blk00000003_sig00000262,
      S => blk00000003_sig00000260,
      O => blk00000003_sig0000025b
    );
  blk00000003_blk000001d3 : XORCY
    port map (
      CI => blk00000003_sig0000025f,
      LI => blk00000003_sig00000260,
      O => blk00000003_sig00000261
    );
  blk00000003_blk000001d2 : MUXCY
    port map (
      CI => blk00000003_sig0000024c,
      DI => blk00000003_sig0000024a,
      S => blk00000003_sig0000024d,
      O => blk00000003_sig0000025e
    );
  blk00000003_blk000001d1 : MUXCY
    port map (
      CI => blk00000003_sig0000025b,
      DI => blk00000003_sig00000245,
      S => blk00000003_sig0000025c,
      O => blk00000003_sig00000258
    );
  blk00000003_blk000001d0 : MUXCY
    port map (
      CI => blk00000003_sig00000258,
      DI => blk00000003_sig00000246,
      S => blk00000003_sig00000259,
      O => blk00000003_sig00000255
    );
  blk00000003_blk000001cf : MUXCY
    port map (
      CI => blk00000003_sig00000255,
      DI => blk00000003_sig00000247,
      S => blk00000003_sig00000256,
      O => blk00000003_sig00000252
    );
  blk00000003_blk000001ce : MUXCY
    port map (
      CI => blk00000003_sig00000252,
      DI => blk00000003_sig00000248,
      S => blk00000003_sig00000253,
      O => blk00000003_sig0000024f
    );
  blk00000003_blk000001cd : MUXCY
    port map (
      CI => blk00000003_sig0000024f,
      DI => blk00000003_sig00000249,
      S => blk00000003_sig00000250,
      O => blk00000003_sig0000024c
    );
  blk00000003_blk000001cc : XORCY
    port map (
      CI => blk00000003_sig0000025b,
      LI => blk00000003_sig0000025c,
      O => blk00000003_sig0000025d
    );
  blk00000003_blk000001cb : XORCY
    port map (
      CI => blk00000003_sig00000258,
      LI => blk00000003_sig00000259,
      O => blk00000003_sig0000025a
    );
  blk00000003_blk000001ca : XORCY
    port map (
      CI => blk00000003_sig00000255,
      LI => blk00000003_sig00000256,
      O => blk00000003_sig00000257
    );
  blk00000003_blk000001c9 : XORCY
    port map (
      CI => blk00000003_sig00000252,
      LI => blk00000003_sig00000253,
      O => blk00000003_sig00000254
    );
  blk00000003_blk000001c8 : XORCY
    port map (
      CI => blk00000003_sig0000024f,
      LI => blk00000003_sig00000250,
      O => blk00000003_sig00000251
    );
  blk00000003_blk000001c7 : XORCY
    port map (
      CI => blk00000003_sig0000024c,
      LI => blk00000003_sig0000024d,
      O => blk00000003_sig0000024e
    );
  blk00000003_blk000001c6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000240,
      Q => blk00000003_sig0000024b
    );
  blk00000003_blk000001c5 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000230,
      Q => blk00000003_sig00000073
    );
  blk00000003_blk000001c4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000233,
      Q => blk00000003_sig0000024a
    );
  blk00000003_blk000001c3 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000236,
      Q => blk00000003_sig00000249
    );
  blk00000003_blk000001c2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000239,
      Q => blk00000003_sig00000248
    );
  blk00000003_blk000001c1 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000023c,
      Q => blk00000003_sig00000247
    );
  blk00000003_blk000001c0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000023f,
      Q => blk00000003_sig00000246
    );
  blk00000003_blk000001bf : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000243,
      Q => blk00000003_sig00000245
    );
  blk00000003_blk000001be : MUXCY
    port map (
      CI => blk00000003_sig00000241,
      DI => blk00000003_sig00000244,
      S => blk00000003_sig00000242,
      O => blk00000003_sig0000023d
    );
  blk00000003_blk000001bd : XORCY
    port map (
      CI => blk00000003_sig00000241,
      LI => blk00000003_sig00000242,
      O => blk00000003_sig00000243
    );
  blk00000003_blk000001bc : MUXCY
    port map (
      CI => blk00000003_sig0000022e,
      DI => blk00000003_sig0000022c,
      S => blk00000003_sig0000022f,
      O => blk00000003_sig00000240
    );
  blk00000003_blk000001bb : MUXCY
    port map (
      CI => blk00000003_sig0000023d,
      DI => blk00000003_sig00000227,
      S => blk00000003_sig0000023e,
      O => blk00000003_sig0000023a
    );
  blk00000003_blk000001ba : MUXCY
    port map (
      CI => blk00000003_sig0000023a,
      DI => blk00000003_sig00000228,
      S => blk00000003_sig0000023b,
      O => blk00000003_sig00000237
    );
  blk00000003_blk000001b9 : MUXCY
    port map (
      CI => blk00000003_sig00000237,
      DI => blk00000003_sig00000229,
      S => blk00000003_sig00000238,
      O => blk00000003_sig00000234
    );
  blk00000003_blk000001b8 : MUXCY
    port map (
      CI => blk00000003_sig00000234,
      DI => blk00000003_sig0000022a,
      S => blk00000003_sig00000235,
      O => blk00000003_sig00000231
    );
  blk00000003_blk000001b7 : MUXCY
    port map (
      CI => blk00000003_sig00000231,
      DI => blk00000003_sig0000022b,
      S => blk00000003_sig00000232,
      O => blk00000003_sig0000022e
    );
  blk00000003_blk000001b6 : XORCY
    port map (
      CI => blk00000003_sig0000023d,
      LI => blk00000003_sig0000023e,
      O => blk00000003_sig0000023f
    );
  blk00000003_blk000001b5 : XORCY
    port map (
      CI => blk00000003_sig0000023a,
      LI => blk00000003_sig0000023b,
      O => blk00000003_sig0000023c
    );
  blk00000003_blk000001b4 : XORCY
    port map (
      CI => blk00000003_sig00000237,
      LI => blk00000003_sig00000238,
      O => blk00000003_sig00000239
    );
  blk00000003_blk000001b3 : XORCY
    port map (
      CI => blk00000003_sig00000234,
      LI => blk00000003_sig00000235,
      O => blk00000003_sig00000236
    );
  blk00000003_blk000001b2 : XORCY
    port map (
      CI => blk00000003_sig00000231,
      LI => blk00000003_sig00000232,
      O => blk00000003_sig00000233
    );
  blk00000003_blk000001b1 : XORCY
    port map (
      CI => blk00000003_sig0000022e,
      LI => blk00000003_sig0000022f,
      O => blk00000003_sig00000230
    );
  blk00000003_blk000001b0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000222,
      Q => blk00000003_sig0000022d
    );
  blk00000003_blk000001af : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000212,
      Q => blk00000003_sig0000007f
    );
  blk00000003_blk000001ae : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000215,
      Q => blk00000003_sig0000022c
    );
  blk00000003_blk000001ad : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000218,
      Q => blk00000003_sig0000022b
    );
  blk00000003_blk000001ac : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000021b,
      Q => blk00000003_sig0000022a
    );
  blk00000003_blk000001ab : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000021e,
      Q => blk00000003_sig00000229
    );
  blk00000003_blk000001aa : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000221,
      Q => blk00000003_sig00000228
    );
  blk00000003_blk000001a9 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000225,
      Q => blk00000003_sig00000227
    );
  blk00000003_blk000001a8 : MUXCY
    port map (
      CI => blk00000003_sig00000223,
      DI => blk00000003_sig00000226,
      S => blk00000003_sig00000224,
      O => blk00000003_sig0000021f
    );
  blk00000003_blk000001a7 : XORCY
    port map (
      CI => blk00000003_sig00000223,
      LI => blk00000003_sig00000224,
      O => blk00000003_sig00000225
    );
  blk00000003_blk000001a6 : MUXCY
    port map (
      CI => blk00000003_sig00000210,
      DI => blk00000003_sig0000020e,
      S => blk00000003_sig00000211,
      O => blk00000003_sig00000222
    );
  blk00000003_blk000001a5 : MUXCY
    port map (
      CI => blk00000003_sig0000021f,
      DI => blk00000003_sig00000209,
      S => blk00000003_sig00000220,
      O => blk00000003_sig0000021c
    );
  blk00000003_blk000001a4 : MUXCY
    port map (
      CI => blk00000003_sig0000021c,
      DI => blk00000003_sig0000020a,
      S => blk00000003_sig0000021d,
      O => blk00000003_sig00000219
    );
  blk00000003_blk000001a3 : MUXCY
    port map (
      CI => blk00000003_sig00000219,
      DI => blk00000003_sig0000020b,
      S => blk00000003_sig0000021a,
      O => blk00000003_sig00000216
    );
  blk00000003_blk000001a2 : MUXCY
    port map (
      CI => blk00000003_sig00000216,
      DI => blk00000003_sig0000020c,
      S => blk00000003_sig00000217,
      O => blk00000003_sig00000213
    );
  blk00000003_blk000001a1 : MUXCY
    port map (
      CI => blk00000003_sig00000213,
      DI => blk00000003_sig0000020d,
      S => blk00000003_sig00000214,
      O => blk00000003_sig00000210
    );
  blk00000003_blk000001a0 : XORCY
    port map (
      CI => blk00000003_sig0000021f,
      LI => blk00000003_sig00000220,
      O => blk00000003_sig00000221
    );
  blk00000003_blk0000019f : XORCY
    port map (
      CI => blk00000003_sig0000021c,
      LI => blk00000003_sig0000021d,
      O => blk00000003_sig0000021e
    );
  blk00000003_blk0000019e : XORCY
    port map (
      CI => blk00000003_sig00000219,
      LI => blk00000003_sig0000021a,
      O => blk00000003_sig0000021b
    );
  blk00000003_blk0000019d : XORCY
    port map (
      CI => blk00000003_sig00000216,
      LI => blk00000003_sig00000217,
      O => blk00000003_sig00000218
    );
  blk00000003_blk0000019c : XORCY
    port map (
      CI => blk00000003_sig00000213,
      LI => blk00000003_sig00000214,
      O => blk00000003_sig00000215
    );
  blk00000003_blk0000019b : XORCY
    port map (
      CI => blk00000003_sig00000210,
      LI => blk00000003_sig00000211,
      O => blk00000003_sig00000212
    );
  blk00000003_blk0000019a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000204,
      Q => blk00000003_sig0000020f
    );
  blk00000003_blk00000199 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001f4,
      Q => blk00000003_sig00000084
    );
  blk00000003_blk00000198 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001f7,
      Q => blk00000003_sig0000020e
    );
  blk00000003_blk00000197 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001fa,
      Q => blk00000003_sig0000020d
    );
  blk00000003_blk00000196 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001fd,
      Q => blk00000003_sig0000020c
    );
  blk00000003_blk00000195 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000200,
      Q => blk00000003_sig0000020b
    );
  blk00000003_blk00000194 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000203,
      Q => blk00000003_sig0000020a
    );
  blk00000003_blk00000193 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000207,
      Q => blk00000003_sig00000209
    );
  blk00000003_blk00000192 : MUXCY
    port map (
      CI => blk00000003_sig00000205,
      DI => blk00000003_sig00000208,
      S => blk00000003_sig00000206,
      O => blk00000003_sig00000201
    );
  blk00000003_blk00000191 : XORCY
    port map (
      CI => blk00000003_sig00000205,
      LI => blk00000003_sig00000206,
      O => blk00000003_sig00000207
    );
  blk00000003_blk00000190 : MUXCY
    port map (
      CI => blk00000003_sig000001f2,
      DI => blk00000003_sig000001f0,
      S => blk00000003_sig000001f3,
      O => blk00000003_sig00000204
    );
  blk00000003_blk0000018f : MUXCY
    port map (
      CI => blk00000003_sig00000201,
      DI => blk00000003_sig000001eb,
      S => blk00000003_sig00000202,
      O => blk00000003_sig000001fe
    );
  blk00000003_blk0000018e : MUXCY
    port map (
      CI => blk00000003_sig000001fe,
      DI => blk00000003_sig000001ec,
      S => blk00000003_sig000001ff,
      O => blk00000003_sig000001fb
    );
  blk00000003_blk0000018d : MUXCY
    port map (
      CI => blk00000003_sig000001fb,
      DI => blk00000003_sig000001ed,
      S => blk00000003_sig000001fc,
      O => blk00000003_sig000001f8
    );
  blk00000003_blk0000018c : MUXCY
    port map (
      CI => blk00000003_sig000001f8,
      DI => blk00000003_sig000001ee,
      S => blk00000003_sig000001f9,
      O => blk00000003_sig000001f5
    );
  blk00000003_blk0000018b : MUXCY
    port map (
      CI => blk00000003_sig000001f5,
      DI => blk00000003_sig000001ef,
      S => blk00000003_sig000001f6,
      O => blk00000003_sig000001f2
    );
  blk00000003_blk0000018a : XORCY
    port map (
      CI => blk00000003_sig00000201,
      LI => blk00000003_sig00000202,
      O => blk00000003_sig00000203
    );
  blk00000003_blk00000189 : XORCY
    port map (
      CI => blk00000003_sig000001fe,
      LI => blk00000003_sig000001ff,
      O => blk00000003_sig00000200
    );
  blk00000003_blk00000188 : XORCY
    port map (
      CI => blk00000003_sig000001fb,
      LI => blk00000003_sig000001fc,
      O => blk00000003_sig000001fd
    );
  blk00000003_blk00000187 : XORCY
    port map (
      CI => blk00000003_sig000001f8,
      LI => blk00000003_sig000001f9,
      O => blk00000003_sig000001fa
    );
  blk00000003_blk00000186 : XORCY
    port map (
      CI => blk00000003_sig000001f5,
      LI => blk00000003_sig000001f6,
      O => blk00000003_sig000001f7
    );
  blk00000003_blk00000185 : XORCY
    port map (
      CI => blk00000003_sig000001f2,
      LI => blk00000003_sig000001f3,
      O => blk00000003_sig000001f4
    );
  blk00000003_blk00000184 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001e6,
      Q => blk00000003_sig000001f1
    );
  blk00000003_blk00000183 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001d6,
      Q => blk00000003_sig00000088
    );
  blk00000003_blk00000182 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001d9,
      Q => blk00000003_sig000001f0
    );
  blk00000003_blk00000181 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001dc,
      Q => blk00000003_sig000001ef
    );
  blk00000003_blk00000180 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001df,
      Q => blk00000003_sig000001ee
    );
  blk00000003_blk0000017f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001e2,
      Q => blk00000003_sig000001ed
    );
  blk00000003_blk0000017e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001e5,
      Q => blk00000003_sig000001ec
    );
  blk00000003_blk0000017d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001e9,
      Q => blk00000003_sig000001eb
    );
  blk00000003_blk0000017c : MUXCY
    port map (
      CI => blk00000003_sig000001e7,
      DI => blk00000003_sig000001ea,
      S => blk00000003_sig000001e8,
      O => blk00000003_sig000001e3
    );
  blk00000003_blk0000017b : XORCY
    port map (
      CI => blk00000003_sig000001e7,
      LI => blk00000003_sig000001e8,
      O => blk00000003_sig000001e9
    );
  blk00000003_blk0000017a : MUXCY
    port map (
      CI => blk00000003_sig000001d4,
      DI => blk00000003_sig000001d2,
      S => blk00000003_sig000001d5,
      O => blk00000003_sig000001e6
    );
  blk00000003_blk00000179 : MUXCY
    port map (
      CI => blk00000003_sig000001e3,
      DI => blk00000003_sig000001cd,
      S => blk00000003_sig000001e4,
      O => blk00000003_sig000001e0
    );
  blk00000003_blk00000178 : MUXCY
    port map (
      CI => blk00000003_sig000001e0,
      DI => blk00000003_sig000001ce,
      S => blk00000003_sig000001e1,
      O => blk00000003_sig000001dd
    );
  blk00000003_blk00000177 : MUXCY
    port map (
      CI => blk00000003_sig000001dd,
      DI => blk00000003_sig000001cf,
      S => blk00000003_sig000001de,
      O => blk00000003_sig000001da
    );
  blk00000003_blk00000176 : MUXCY
    port map (
      CI => blk00000003_sig000001da,
      DI => blk00000003_sig000001d0,
      S => blk00000003_sig000001db,
      O => blk00000003_sig000001d7
    );
  blk00000003_blk00000175 : MUXCY
    port map (
      CI => blk00000003_sig000001d7,
      DI => blk00000003_sig000001d1,
      S => blk00000003_sig000001d8,
      O => blk00000003_sig000001d4
    );
  blk00000003_blk00000174 : XORCY
    port map (
      CI => blk00000003_sig000001e3,
      LI => blk00000003_sig000001e4,
      O => blk00000003_sig000001e5
    );
  blk00000003_blk00000173 : XORCY
    port map (
      CI => blk00000003_sig000001e0,
      LI => blk00000003_sig000001e1,
      O => blk00000003_sig000001e2
    );
  blk00000003_blk00000172 : XORCY
    port map (
      CI => blk00000003_sig000001dd,
      LI => blk00000003_sig000001de,
      O => blk00000003_sig000001df
    );
  blk00000003_blk00000171 : XORCY
    port map (
      CI => blk00000003_sig000001da,
      LI => blk00000003_sig000001db,
      O => blk00000003_sig000001dc
    );
  blk00000003_blk00000170 : XORCY
    port map (
      CI => blk00000003_sig000001d7,
      LI => blk00000003_sig000001d8,
      O => blk00000003_sig000001d9
    );
  blk00000003_blk0000016f : XORCY
    port map (
      CI => blk00000003_sig000001d4,
      LI => blk00000003_sig000001d5,
      O => blk00000003_sig000001d6
    );
  blk00000003_blk0000016e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001c8,
      Q => blk00000003_sig000001d3
    );
  blk00000003_blk0000016d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001b8,
      Q => blk00000003_sig0000008b
    );
  blk00000003_blk0000016c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001bb,
      Q => blk00000003_sig000001d2
    );
  blk00000003_blk0000016b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001be,
      Q => blk00000003_sig000001d1
    );
  blk00000003_blk0000016a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001c1,
      Q => blk00000003_sig000001d0
    );
  blk00000003_blk00000169 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001c4,
      Q => blk00000003_sig000001cf
    );
  blk00000003_blk00000168 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001c7,
      Q => blk00000003_sig000001ce
    );
  blk00000003_blk00000167 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001cb,
      Q => blk00000003_sig000001cd
    );
  blk00000003_blk00000166 : MUXCY
    port map (
      CI => blk00000003_sig000001c9,
      DI => blk00000003_sig000001cc,
      S => blk00000003_sig000001ca,
      O => blk00000003_sig000001c5
    );
  blk00000003_blk00000165 : XORCY
    port map (
      CI => blk00000003_sig000001c9,
      LI => blk00000003_sig000001ca,
      O => blk00000003_sig000001cb
    );
  blk00000003_blk00000164 : MUXCY
    port map (
      CI => blk00000003_sig000001b6,
      DI => blk00000003_sig000001b5,
      S => blk00000003_sig000001b7,
      O => blk00000003_sig000001c8
    );
  blk00000003_blk00000163 : MUXCY
    port map (
      CI => blk00000003_sig000001c5,
      DI => blk00000003_sig000001b0,
      S => blk00000003_sig000001c6,
      O => blk00000003_sig000001c2
    );
  blk00000003_blk00000162 : MUXCY
    port map (
      CI => blk00000003_sig000001c2,
      DI => blk00000003_sig000001b1,
      S => blk00000003_sig000001c3,
      O => blk00000003_sig000001bf
    );
  blk00000003_blk00000161 : MUXCY
    port map (
      CI => blk00000003_sig000001bf,
      DI => blk00000003_sig000001b2,
      S => blk00000003_sig000001c0,
      O => blk00000003_sig000001bc
    );
  blk00000003_blk00000160 : MUXCY
    port map (
      CI => blk00000003_sig000001bc,
      DI => blk00000003_sig000001b3,
      S => blk00000003_sig000001bd,
      O => blk00000003_sig000001b9
    );
  blk00000003_blk0000015f : MUXCY
    port map (
      CI => blk00000003_sig000001b9,
      DI => blk00000003_sig000001b4,
      S => blk00000003_sig000001ba,
      O => blk00000003_sig000001b6
    );
  blk00000003_blk0000015e : XORCY
    port map (
      CI => blk00000003_sig000001c5,
      LI => blk00000003_sig000001c6,
      O => blk00000003_sig000001c7
    );
  blk00000003_blk0000015d : XORCY
    port map (
      CI => blk00000003_sig000001c2,
      LI => blk00000003_sig000001c3,
      O => blk00000003_sig000001c4
    );
  blk00000003_blk0000015c : XORCY
    port map (
      CI => blk00000003_sig000001bf,
      LI => blk00000003_sig000001c0,
      O => blk00000003_sig000001c1
    );
  blk00000003_blk0000015b : XORCY
    port map (
      CI => blk00000003_sig000001bc,
      LI => blk00000003_sig000001bd,
      O => blk00000003_sig000001be
    );
  blk00000003_blk0000015a : XORCY
    port map (
      CI => blk00000003_sig000001b9,
      LI => blk00000003_sig000001ba,
      O => blk00000003_sig000001bb
    );
  blk00000003_blk00000159 : XORCY
    port map (
      CI => blk00000003_sig000001b6,
      LI => blk00000003_sig000001b7,
      O => blk00000003_sig000001b8
    );
  blk00000003_blk00000158 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000019e,
      Q => blk00000003_sig0000008d
    );
  blk00000003_blk00000157 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001a1,
      Q => blk00000003_sig000001b5
    );
  blk00000003_blk00000156 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001a4,
      Q => blk00000003_sig000001b4
    );
  blk00000003_blk00000155 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001a7,
      Q => blk00000003_sig000001b3
    );
  blk00000003_blk00000154 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001aa,
      Q => blk00000003_sig000001b2
    );
  blk00000003_blk00000153 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001ad,
      Q => blk00000003_sig000001b1
    );
  blk00000003_blk00000152 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000001af,
      Q => blk00000003_sig000001b0
    );
  blk00000003_blk00000151 : MUXCY
    port map (
      CI => NlwRenamedSig_OI_rfd,
      DI => blk00000003_sig0000017d,
      S => blk00000003_sig000001ae,
      O => blk00000003_sig000001ab
    );
  blk00000003_blk00000150 : XORCY
    port map (
      CI => NlwRenamedSig_OI_rfd,
      LI => blk00000003_sig000001ae,
      O => blk00000003_sig000001af
    );
  blk00000003_blk0000014f : MUXCY
    port map (
      CI => blk00000003_sig0000019d,
      DI => blk00000003_sig0000004f,
      S => NlwRenamedSig_OI_rfd,
      O => NLW_blk00000003_blk0000014f_O_UNCONNECTED
    );
  blk00000003_blk0000014e : MUXCY
    port map (
      CI => blk00000003_sig000001ab,
      DI => blk00000003_sig0000004f,
      S => blk00000003_sig000001ac,
      O => blk00000003_sig000001a8
    );
  blk00000003_blk0000014d : MUXCY
    port map (
      CI => blk00000003_sig000001a8,
      DI => blk00000003_sig0000004f,
      S => blk00000003_sig000001a9,
      O => blk00000003_sig000001a5
    );
  blk00000003_blk0000014c : MUXCY
    port map (
      CI => blk00000003_sig000001a5,
      DI => blk00000003_sig0000004f,
      S => blk00000003_sig000001a6,
      O => blk00000003_sig000001a2
    );
  blk00000003_blk0000014b : MUXCY
    port map (
      CI => blk00000003_sig000001a2,
      DI => blk00000003_sig0000004f,
      S => blk00000003_sig000001a3,
      O => blk00000003_sig0000019f
    );
  blk00000003_blk0000014a : MUXCY
    port map (
      CI => blk00000003_sig0000019f,
      DI => blk00000003_sig0000004f,
      S => blk00000003_sig000001a0,
      O => blk00000003_sig0000019d
    );
  blk00000003_blk00000149 : XORCY
    port map (
      CI => blk00000003_sig000001ab,
      LI => blk00000003_sig000001ac,
      O => blk00000003_sig000001ad
    );
  blk00000003_blk00000148 : XORCY
    port map (
      CI => blk00000003_sig000001a8,
      LI => blk00000003_sig000001a9,
      O => blk00000003_sig000001aa
    );
  blk00000003_blk00000147 : XORCY
    port map (
      CI => blk00000003_sig000001a5,
      LI => blk00000003_sig000001a6,
      O => blk00000003_sig000001a7
    );
  blk00000003_blk00000146 : XORCY
    port map (
      CI => blk00000003_sig000001a2,
      LI => blk00000003_sig000001a3,
      O => blk00000003_sig000001a4
    );
  blk00000003_blk00000145 : XORCY
    port map (
      CI => blk00000003_sig0000019f,
      LI => blk00000003_sig000001a0,
      O => blk00000003_sig000001a1
    );
  blk00000003_blk00000144 : XORCY
    port map (
      CI => blk00000003_sig0000019d,
      LI => NlwRenamedSig_OI_rfd,
      O => blk00000003_sig0000019e
    );
  blk00000003_blk00000143 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(0),
      Q => blk00000003_sig0000019c
    );
  blk00000003_blk00000142 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(1),
      Q => blk00000003_sig0000019b
    );
  blk00000003_blk00000141 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(2),
      Q => blk00000003_sig0000019a
    );
  blk00000003_blk00000140 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(3),
      Q => blk00000003_sig00000199
    );
  blk00000003_blk0000013f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(4),
      Q => blk00000003_sig00000198
    );
  blk00000003_blk0000013e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(5),
      Q => blk00000003_sig00000197
    );
  blk00000003_blk0000013d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(6),
      Q => blk00000003_sig00000196
    );
  blk00000003_blk0000013c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(7),
      Q => blk00000003_sig00000195
    );
  blk00000003_blk0000013b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(8),
      Q => blk00000003_sig00000194
    );
  blk00000003_blk0000013a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(9),
      Q => blk00000003_sig00000193
    );
  blk00000003_blk00000139 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(10),
      Q => blk00000003_sig00000192
    );
  blk00000003_blk00000138 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(11),
      Q => blk00000003_sig00000191
    );
  blk00000003_blk00000137 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(12),
      Q => blk00000003_sig00000190
    );
  blk00000003_blk00000136 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(13),
      Q => blk00000003_sig0000018f
    );
  blk00000003_blk00000135 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(14),
      Q => blk00000003_sig0000018e
    );
  blk00000003_blk00000134 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(15),
      Q => blk00000003_sig0000018d
    );
  blk00000003_blk00000133 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(16),
      Q => blk00000003_sig0000018c
    );
  blk00000003_blk00000132 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(17),
      Q => blk00000003_sig0000018b
    );
  blk00000003_blk00000131 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(18),
      Q => blk00000003_sig0000018a
    );
  blk00000003_blk00000130 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(19),
      Q => blk00000003_sig00000189
    );
  blk00000003_blk0000012f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(20),
      Q => blk00000003_sig00000188
    );
  blk00000003_blk0000012e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(21),
      Q => blk00000003_sig00000187
    );
  blk00000003_blk0000012d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(22),
      Q => blk00000003_sig00000186
    );
  blk00000003_blk0000012c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(23),
      Q => blk00000003_sig00000185
    );
  blk00000003_blk0000012b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(24),
      Q => blk00000003_sig00000184
    );
  blk00000003_blk0000012a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(25),
      Q => blk00000003_sig00000183
    );
  blk00000003_blk00000129 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(26),
      Q => blk00000003_sig00000182
    );
  blk00000003_blk00000128 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(27),
      Q => blk00000003_sig00000181
    );
  blk00000003_blk00000127 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(28),
      Q => blk00000003_sig00000180
    );
  blk00000003_blk00000126 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(29),
      Q => blk00000003_sig0000017f
    );
  blk00000003_blk00000125 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(30),
      Q => blk00000003_sig0000017e
    );
  blk00000003_blk00000124 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => dividend(31),
      Q => blk00000003_sig0000017d
    );
  blk00000003_blk00000123 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000017c,
      Q => quotient(0)
    );
  blk00000003_blk00000122 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000017b,
      Q => quotient(1)
    );
  blk00000003_blk00000121 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000017a,
      Q => quotient(2)
    );
  blk00000003_blk00000120 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000179,
      Q => quotient(3)
    );
  blk00000003_blk0000011f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000178,
      Q => quotient(4)
    );
  blk00000003_blk0000011e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000177,
      Q => quotient(5)
    );
  blk00000003_blk0000011d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000176,
      Q => quotient(6)
    );
  blk00000003_blk0000011c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000175,
      Q => quotient(7)
    );
  blk00000003_blk0000011b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000174,
      Q => quotient(8)
    );
  blk00000003_blk0000011a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000173,
      Q => quotient(9)
    );
  blk00000003_blk00000119 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000172,
      Q => quotient(10)
    );
  blk00000003_blk00000118 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000171,
      Q => quotient(11)
    );
  blk00000003_blk00000117 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000170,
      Q => quotient(12)
    );
  blk00000003_blk00000116 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000016f,
      Q => quotient(13)
    );
  blk00000003_blk00000115 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000016e,
      Q => quotient(14)
    );
  blk00000003_blk00000114 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000016d,
      Q => quotient(15)
    );
  blk00000003_blk00000113 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000016c,
      Q => quotient(16)
    );
  blk00000003_blk00000112 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000016b,
      Q => quotient(17)
    );
  blk00000003_blk00000111 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000016a,
      Q => quotient(18)
    );
  blk00000003_blk00000110 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000169,
      Q => quotient(19)
    );
  blk00000003_blk0000010f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000168,
      Q => quotient(20)
    );
  blk00000003_blk0000010e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000167,
      Q => quotient(21)
    );
  blk00000003_blk0000010d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000166,
      Q => quotient(22)
    );
  blk00000003_blk0000010c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000165,
      Q => quotient(23)
    );
  blk00000003_blk0000010b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000164,
      Q => quotient(24)
    );
  blk00000003_blk0000010a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000163,
      Q => quotient(25)
    );
  blk00000003_blk00000109 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000162,
      Q => quotient(26)
    );
  blk00000003_blk00000108 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000161,
      Q => quotient(27)
    );
  blk00000003_blk00000107 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000160,
      Q => quotient(28)
    );
  blk00000003_blk00000106 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000015f,
      Q => quotient(29)
    );
  blk00000003_blk00000105 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000015e,
      Q => quotient(30)
    );
  blk00000003_blk00000104 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000015d,
      Q => quotient(31)
    );
  blk00000003_blk00000103 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000156,
      Q => blk00000003_sig0000015c
    );
  blk00000003_blk00000102 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000155,
      Q => blk00000003_sig0000015b
    );
  blk00000003_blk00000101 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000154,
      Q => blk00000003_sig0000015a
    );
  blk00000003_blk00000100 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000153,
      Q => blk00000003_sig00000159
    );
  blk00000003_blk000000ff : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000152,
      Q => blk00000003_sig00000158
    );
  blk00000003_blk000000fe : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000151,
      Q => blk00000003_sig00000157
    );
  blk00000003_blk000000fd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000150,
      Q => blk00000003_sig00000156
    );
  blk00000003_blk000000fc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000014f,
      Q => blk00000003_sig00000155
    );
  blk00000003_blk000000fb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000014e,
      Q => blk00000003_sig00000154
    );
  blk00000003_blk000000fa : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000014d,
      Q => blk00000003_sig00000153
    );
  blk00000003_blk000000f9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000014c,
      Q => blk00000003_sig00000152
    );
  blk00000003_blk000000f8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000014b,
      Q => blk00000003_sig00000151
    );
  blk00000003_blk000000f7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000014a,
      Q => blk00000003_sig00000150
    );
  blk00000003_blk000000f6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000149,
      Q => blk00000003_sig0000014f
    );
  blk00000003_blk000000f5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000148,
      Q => blk00000003_sig0000014e
    );
  blk00000003_blk000000f4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000147,
      Q => blk00000003_sig0000014d
    );
  blk00000003_blk000000f3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000146,
      Q => blk00000003_sig0000014c
    );
  blk00000003_blk000000f2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000145,
      Q => blk00000003_sig0000014b
    );
  blk00000003_blk000000f1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000144,
      Q => blk00000003_sig0000014a
    );
  blk00000003_blk000000f0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000143,
      Q => blk00000003_sig00000149
    );
  blk00000003_blk000000ef : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000142,
      Q => blk00000003_sig00000148
    );
  blk00000003_blk000000ee : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000141,
      Q => blk00000003_sig00000147
    );
  blk00000003_blk000000ed : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000140,
      Q => blk00000003_sig00000146
    );
  blk00000003_blk000000ec : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000013f,
      Q => blk00000003_sig00000145
    );
  blk00000003_blk000000eb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000013e,
      Q => blk00000003_sig00000144
    );
  blk00000003_blk000000ea : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000013d,
      Q => blk00000003_sig00000143
    );
  blk00000003_blk000000e9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000013c,
      Q => blk00000003_sig00000142
    );
  blk00000003_blk000000e8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000013b,
      Q => blk00000003_sig00000141
    );
  blk00000003_blk000000e7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000013a,
      Q => blk00000003_sig00000140
    );
  blk00000003_blk000000e6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000139,
      Q => blk00000003_sig0000013f
    );
  blk00000003_blk000000e5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000138,
      Q => blk00000003_sig0000013e
    );
  blk00000003_blk000000e4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000137,
      Q => blk00000003_sig0000013d
    );
  blk00000003_blk000000e3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000136,
      Q => blk00000003_sig0000013c
    );
  blk00000003_blk000000e2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000135,
      Q => blk00000003_sig0000013b
    );
  blk00000003_blk000000e1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000134,
      Q => blk00000003_sig0000013a
    );
  blk00000003_blk000000e0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000133,
      Q => blk00000003_sig00000139
    );
  blk00000003_blk000000df : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000132,
      Q => blk00000003_sig00000138
    );
  blk00000003_blk000000de : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000131,
      Q => blk00000003_sig00000137
    );
  blk00000003_blk000000dd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000130,
      Q => blk00000003_sig00000136
    );
  blk00000003_blk000000dc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000012f,
      Q => blk00000003_sig00000135
    );
  blk00000003_blk000000db : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000012e,
      Q => blk00000003_sig00000134
    );
  blk00000003_blk000000da : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000012d,
      Q => blk00000003_sig00000133
    );
  blk00000003_blk000000d9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000012c,
      Q => blk00000003_sig00000132
    );
  blk00000003_blk000000d8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000012b,
      Q => blk00000003_sig00000131
    );
  blk00000003_blk000000d7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000012a,
      Q => blk00000003_sig00000130
    );
  blk00000003_blk000000d6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000129,
      Q => blk00000003_sig0000012f
    );
  blk00000003_blk000000d5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000128,
      Q => blk00000003_sig0000012e
    );
  blk00000003_blk000000d4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000127,
      Q => blk00000003_sig0000012d
    );
  blk00000003_blk000000d3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000126,
      Q => blk00000003_sig0000012c
    );
  blk00000003_blk000000d2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000125,
      Q => blk00000003_sig0000012b
    );
  blk00000003_blk000000d1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000124,
      Q => blk00000003_sig0000012a
    );
  blk00000003_blk000000d0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000123,
      Q => blk00000003_sig00000129
    );
  blk00000003_blk000000cf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000122,
      Q => blk00000003_sig00000128
    );
  blk00000003_blk000000ce : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000121,
      Q => blk00000003_sig00000127
    );
  blk00000003_blk000000cd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000120,
      Q => blk00000003_sig00000126
    );
  blk00000003_blk000000cc : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000011f,
      Q => blk00000003_sig00000125
    );
  blk00000003_blk000000cb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000011e,
      Q => blk00000003_sig00000124
    );
  blk00000003_blk000000ca : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000011d,
      Q => blk00000003_sig00000123
    );
  blk00000003_blk000000c9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000011c,
      Q => blk00000003_sig00000122
    );
  blk00000003_blk000000c8 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000011b,
      Q => blk00000003_sig00000121
    );
  blk00000003_blk000000c7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000011a,
      Q => blk00000003_sig00000120
    );
  blk00000003_blk000000c6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000119,
      Q => blk00000003_sig0000011f
    );
  blk00000003_blk000000c5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000118,
      Q => blk00000003_sig0000011e
    );
  blk00000003_blk000000c4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000117,
      Q => blk00000003_sig0000011d
    );
  blk00000003_blk000000c3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000116,
      Q => blk00000003_sig0000011c
    );
  blk00000003_blk000000c2 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000115,
      Q => blk00000003_sig0000011b
    );
  blk00000003_blk000000c1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000114,
      Q => blk00000003_sig0000011a
    );
  blk00000003_blk000000c0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000113,
      Q => blk00000003_sig00000119
    );
  blk00000003_blk000000bf : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000112,
      Q => blk00000003_sig00000118
    );
  blk00000003_blk000000be : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000111,
      Q => blk00000003_sig00000117
    );
  blk00000003_blk000000bd : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000110,
      Q => blk00000003_sig00000116
    );
  blk00000003_blk000000bc : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000010f,
      Q => blk00000003_sig00000115
    );
  blk00000003_blk000000bb : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000010e,
      Q => blk00000003_sig00000114
    );
  blk00000003_blk000000ba : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000010d,
      Q => blk00000003_sig00000113
    );
  blk00000003_blk000000b9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000010c,
      Q => blk00000003_sig00000112
    );
  blk00000003_blk000000b8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000010b,
      Q => blk00000003_sig00000111
    );
  blk00000003_blk000000b7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000010a,
      Q => blk00000003_sig00000110
    );
  blk00000003_blk000000b6 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000109,
      Q => blk00000003_sig0000010f
    );
  blk00000003_blk000000b5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000108,
      Q => blk00000003_sig0000010e
    );
  blk00000003_blk000000b4 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000107,
      Q => blk00000003_sig0000010d
    );
  blk00000003_blk000000b3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000106,
      Q => blk00000003_sig0000010c
    );
  blk00000003_blk000000b2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000105,
      Q => blk00000003_sig0000010b
    );
  blk00000003_blk000000b1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000104,
      Q => blk00000003_sig0000010a
    );
  blk00000003_blk000000b0 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000103,
      Q => blk00000003_sig00000109
    );
  blk00000003_blk000000af : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000102,
      Q => blk00000003_sig00000108
    );
  blk00000003_blk000000ae : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000101,
      Q => blk00000003_sig00000107
    );
  blk00000003_blk000000ad : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000100,
      Q => blk00000003_sig00000106
    );
  blk00000003_blk000000ac : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ff,
      Q => blk00000003_sig00000105
    );
  blk00000003_blk000000ab : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000fe,
      Q => blk00000003_sig00000104
    );
  blk00000003_blk000000aa : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000fd,
      Q => blk00000003_sig00000103
    );
  blk00000003_blk000000a9 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000fc,
      Q => blk00000003_sig00000102
    );
  blk00000003_blk000000a8 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000fb,
      Q => blk00000003_sig00000101
    );
  blk00000003_blk000000a7 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000fa,
      Q => blk00000003_sig00000100
    );
  blk00000003_blk000000a6 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f9,
      Q => blk00000003_sig000000ff
    );
  blk00000003_blk000000a5 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f8,
      Q => blk00000003_sig000000fe
    );
  blk00000003_blk000000a4 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f7,
      Q => blk00000003_sig000000fd
    );
  blk00000003_blk000000a3 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f6,
      Q => blk00000003_sig000000fc
    );
  blk00000003_blk000000a2 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f5,
      Q => blk00000003_sig000000fb
    );
  blk00000003_blk000000a1 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f4,
      Q => blk00000003_sig000000fa
    );
  blk00000003_blk000000a0 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f3,
      Q => blk00000003_sig000000f9
    );
  blk00000003_blk0000009f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f2,
      Q => blk00000003_sig000000f8
    );
  blk00000003_blk0000009e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f1,
      Q => blk00000003_sig000000f7
    );
  blk00000003_blk0000009d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000f0,
      Q => blk00000003_sig000000f6
    );
  blk00000003_blk0000009c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ef,
      Q => blk00000003_sig000000f5
    );
  blk00000003_blk0000009b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ee,
      Q => blk00000003_sig000000f4
    );
  blk00000003_blk0000009a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ed,
      Q => blk00000003_sig000000f3
    );
  blk00000003_blk00000099 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ec,
      Q => blk00000003_sig000000f2
    );
  blk00000003_blk00000098 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000eb,
      Q => blk00000003_sig000000f1
    );
  blk00000003_blk00000097 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ea,
      Q => blk00000003_sig000000f0
    );
  blk00000003_blk00000096 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e9,
      Q => blk00000003_sig000000ef
    );
  blk00000003_blk00000095 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e8,
      Q => blk00000003_sig000000ee
    );
  blk00000003_blk00000094 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e7,
      Q => blk00000003_sig000000ed
    );
  blk00000003_blk00000093 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e6,
      Q => blk00000003_sig000000ec
    );
  blk00000003_blk00000092 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e5,
      Q => blk00000003_sig000000eb
    );
  blk00000003_blk00000091 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e4,
      Q => blk00000003_sig000000ea
    );
  blk00000003_blk00000090 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e3,
      Q => blk00000003_sig000000e9
    );
  blk00000003_blk0000008f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e2,
      Q => blk00000003_sig000000e8
    );
  blk00000003_blk0000008e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e1,
      Q => blk00000003_sig000000e7
    );
  blk00000003_blk0000008d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000e0,
      Q => blk00000003_sig000000e6
    );
  blk00000003_blk0000008c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000df,
      Q => blk00000003_sig000000e5
    );
  blk00000003_blk0000008b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000de,
      Q => blk00000003_sig000000e4
    );
  blk00000003_blk0000008a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000dd,
      Q => blk00000003_sig000000e3
    );
  blk00000003_blk00000089 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000dc,
      Q => blk00000003_sig000000e2
    );
  blk00000003_blk00000088 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000db,
      Q => blk00000003_sig000000e1
    );
  blk00000003_blk00000087 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000da,
      Q => blk00000003_sig000000e0
    );
  blk00000003_blk00000086 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d9,
      Q => blk00000003_sig000000df
    );
  blk00000003_blk00000085 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d8,
      Q => blk00000003_sig000000de
    );
  blk00000003_blk00000084 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d7,
      Q => blk00000003_sig000000dd
    );
  blk00000003_blk00000083 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d6,
      Q => blk00000003_sig000000dc
    );
  blk00000003_blk00000082 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d5,
      Q => blk00000003_sig000000db
    );
  blk00000003_blk00000081 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d4,
      Q => blk00000003_sig000000da
    );
  blk00000003_blk00000080 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d3,
      Q => blk00000003_sig000000d9
    );
  blk00000003_blk0000007f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d2,
      Q => blk00000003_sig000000d8
    );
  blk00000003_blk0000007e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d1,
      Q => blk00000003_sig000000d7
    );
  blk00000003_blk0000007d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000d0,
      Q => blk00000003_sig000000d6
    );
  blk00000003_blk0000007c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000cf,
      Q => blk00000003_sig000000d5
    );
  blk00000003_blk0000007b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ce,
      Q => blk00000003_sig000000d4
    );
  blk00000003_blk0000007a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000cd,
      Q => blk00000003_sig000000d3
    );
  blk00000003_blk00000079 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000cc,
      Q => blk00000003_sig000000d2
    );
  blk00000003_blk00000078 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000cb,
      Q => blk00000003_sig000000d1
    );
  blk00000003_blk00000077 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ca,
      Q => blk00000003_sig000000d0
    );
  blk00000003_blk00000076 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c9,
      Q => blk00000003_sig000000cf
    );
  blk00000003_blk00000075 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c8,
      Q => blk00000003_sig000000ce
    );
  blk00000003_blk00000074 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c7,
      Q => blk00000003_sig000000cd
    );
  blk00000003_blk00000073 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c6,
      Q => blk00000003_sig000000cc
    );
  blk00000003_blk00000072 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c5,
      Q => blk00000003_sig000000cb
    );
  blk00000003_blk00000071 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c4,
      Q => blk00000003_sig000000ca
    );
  blk00000003_blk00000070 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c3,
      Q => blk00000003_sig000000c9
    );
  blk00000003_blk0000006f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c2,
      Q => blk00000003_sig000000c8
    );
  blk00000003_blk0000006e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c1,
      Q => blk00000003_sig000000c7
    );
  blk00000003_blk0000006d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000c0,
      Q => blk00000003_sig000000c6
    );
  blk00000003_blk0000006c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000bf,
      Q => blk00000003_sig000000c5
    );
  blk00000003_blk0000006b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000be,
      Q => blk00000003_sig000000c4
    );
  blk00000003_blk0000006a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000bd,
      Q => blk00000003_sig000000c3
    );
  blk00000003_blk00000069 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000bc,
      Q => blk00000003_sig000000c2
    );
  blk00000003_blk00000068 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000bb,
      Q => blk00000003_sig000000c1
    );
  blk00000003_blk00000067 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ba,
      Q => blk00000003_sig000000c0
    );
  blk00000003_blk00000066 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b9,
      Q => blk00000003_sig000000bf
    );
  blk00000003_blk00000065 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b8,
      Q => blk00000003_sig000000be
    );
  blk00000003_blk00000064 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b7,
      Q => blk00000003_sig000000bd
    );
  blk00000003_blk00000063 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b6,
      Q => blk00000003_sig000000bc
    );
  blk00000003_blk00000062 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b5,
      Q => blk00000003_sig000000bb
    );
  blk00000003_blk00000061 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b4,
      Q => blk00000003_sig000000ba
    );
  blk00000003_blk00000060 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b3,
      Q => blk00000003_sig000000b9
    );
  blk00000003_blk0000005f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b2,
      Q => blk00000003_sig000000b8
    );
  blk00000003_blk0000005e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b1,
      Q => blk00000003_sig000000b7
    );
  blk00000003_blk0000005d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000b0,
      Q => blk00000003_sig000000b6
    );
  blk00000003_blk0000005c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000af,
      Q => blk00000003_sig000000b5
    );
  blk00000003_blk0000005b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ae,
      Q => blk00000003_sig000000b4
    );
  blk00000003_blk0000005a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ad,
      Q => blk00000003_sig000000b3
    );
  blk00000003_blk00000059 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ac,
      Q => blk00000003_sig000000b2
    );
  blk00000003_blk00000058 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000ab,
      Q => blk00000003_sig000000b1
    );
  blk00000003_blk00000057 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000aa,
      Q => blk00000003_sig000000b0
    );
  blk00000003_blk00000056 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a9,
      Q => blk00000003_sig000000af
    );
  blk00000003_blk00000055 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a8,
      Q => blk00000003_sig000000ae
    );
  blk00000003_blk00000054 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a7,
      Q => blk00000003_sig000000ad
    );
  blk00000003_blk00000053 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a6,
      Q => blk00000003_sig000000ac
    );
  blk00000003_blk00000052 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a5,
      Q => blk00000003_sig000000ab
    );
  blk00000003_blk00000051 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a4,
      Q => blk00000003_sig000000aa
    );
  blk00000003_blk00000050 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a3,
      Q => blk00000003_sig000000a9
    );
  blk00000003_blk0000004f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a2,
      Q => blk00000003_sig000000a8
    );
  blk00000003_blk0000004e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a1,
      Q => blk00000003_sig000000a7
    );
  blk00000003_blk0000004d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig000000a0,
      Q => blk00000003_sig000000a6
    );
  blk00000003_blk0000004c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000009f,
      Q => blk00000003_sig000000a5
    );
  blk00000003_blk0000004b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000009e,
      Q => blk00000003_sig000000a4
    );
  blk00000003_blk0000004a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000009d,
      Q => blk00000003_sig000000a3
    );
  blk00000003_blk00000049 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000009c,
      Q => blk00000003_sig000000a2
    );
  blk00000003_blk00000048 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000009b,
      Q => blk00000003_sig000000a1
    );
  blk00000003_blk00000047 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000009a,
      Q => blk00000003_sig000000a0
    );
  blk00000003_blk00000046 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000099,
      Q => blk00000003_sig0000009f
    );
  blk00000003_blk00000045 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000098,
      Q => blk00000003_sig0000009e
    );
  blk00000003_blk00000044 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000097,
      Q => blk00000003_sig0000009d
    );
  blk00000003_blk00000043 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(5),
      Q => blk00000003_sig0000009c
    );
  blk00000003_blk00000042 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(4),
      Q => blk00000003_sig0000009b
    );
  blk00000003_blk00000041 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(3),
      Q => blk00000003_sig0000009a
    );
  blk00000003_blk00000040 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(2),
      Q => blk00000003_sig00000099
    );
  blk00000003_blk0000003f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(1),
      Q => blk00000003_sig00000098
    );
  blk00000003_blk0000003e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => divisor(0),
      Q => blk00000003_sig00000097
    );
  blk00000003_blk0000003d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000052,
      Q => blk00000003_sig00000096
    );
  blk00000003_blk0000003c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007e,
      Q => blk00000003_sig00000095
    );
  blk00000003_blk0000003b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007c,
      Q => blk00000003_sig00000094
    );
  blk00000003_blk0000003a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007a,
      Q => blk00000003_sig00000093
    );
  blk00000003_blk00000039 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000078,
      Q => blk00000003_sig00000092
    );
  blk00000003_blk00000038 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000076,
      Q => blk00000003_sig00000091
    );
  blk00000003_blk00000037 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000074,
      Q => blk00000003_sig00000090
    );
  blk00000003_blk00000036 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000008e,
      Q => blk00000003_sig0000008f
    );
  blk00000003_blk00000035 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000008d,
      Q => blk00000003_sig0000008c
    );
  blk00000003_blk00000034 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000008c,
      Q => blk00000003_sig0000008a
    );
  blk00000003_blk00000033 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000008b,
      Q => blk00000003_sig00000089
    );
  blk00000003_blk00000032 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000008a,
      Q => blk00000003_sig00000087
    );
  blk00000003_blk00000031 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000089,
      Q => blk00000003_sig00000086
    );
  blk00000003_blk00000030 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000088,
      Q => blk00000003_sig00000085
    );
  blk00000003_blk0000002f : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000087,
      Q => blk00000003_sig00000083
    );
  blk00000003_blk0000002e : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000086,
      Q => blk00000003_sig00000082
    );
  blk00000003_blk0000002d : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000085,
      Q => blk00000003_sig00000081
    );
  blk00000003_blk0000002c : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000084,
      Q => blk00000003_sig00000080
    );
  blk00000003_blk0000002b : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000083,
      Q => blk00000003_sig0000007d
    );
  blk00000003_blk0000002a : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000082,
      Q => blk00000003_sig0000007b
    );
  blk00000003_blk00000029 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000081,
      Q => blk00000003_sig00000079
    );
  blk00000003_blk00000028 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000080,
      Q => blk00000003_sig00000077
    );
  blk00000003_blk00000027 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007f,
      Q => blk00000003_sig00000075
    );
  blk00000003_blk00000026 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007d,
      Q => blk00000003_sig0000007e
    );
  blk00000003_blk00000025 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000007b,
      Q => blk00000003_sig0000007c
    );
  blk00000003_blk00000024 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000079,
      Q => blk00000003_sig0000007a
    );
  blk00000003_blk00000023 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000077,
      Q => blk00000003_sig00000078
    );
  blk00000003_blk00000022 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000075,
      Q => blk00000003_sig00000076
    );
  blk00000003_blk00000021 : FDE
    generic map(
      INIT => '1'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000073,
      Q => blk00000003_sig00000074
    );
  blk00000003_blk00000020 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000071,
      Q => blk00000003_sig00000072
    );
  blk00000003_blk0000001f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000070,
      Q => blk00000003_sig00000069
    );
  blk00000003_blk0000001e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006f,
      Q => blk00000003_sig00000068
    );
  blk00000003_blk0000001d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006e,
      Q => blk00000003_sig00000067
    );
  blk00000003_blk0000001c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006d,
      Q => blk00000003_sig00000066
    );
  blk00000003_blk0000001b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006c,
      Q => blk00000003_sig00000065
    );
  blk00000003_blk0000001a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000006b,
      Q => blk00000003_sig00000064
    );
  blk00000003_blk00000019 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000069,
      Q => blk00000003_sig0000006a
    );
  blk00000003_blk00000018 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000068,
      Q => blk00000003_sig00000062
    );
  blk00000003_blk00000017 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000067,
      Q => blk00000003_sig00000061
    );
  blk00000003_blk00000016 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000066,
      Q => blk00000003_sig00000060
    );
  blk00000003_blk00000015 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000065,
      Q => blk00000003_sig0000005f
    );
  blk00000003_blk00000014 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000064,
      Q => blk00000003_sig0000005e
    );
  blk00000003_blk00000013 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000062,
      Q => blk00000003_sig00000063
    );
  blk00000003_blk00000012 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000061,
      Q => blk00000003_sig0000005c
    );
  blk00000003_blk00000011 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000060,
      Q => blk00000003_sig0000005b
    );
  blk00000003_blk00000010 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000005f,
      Q => blk00000003_sig0000005a
    );
  blk00000003_blk0000000f : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000005e,
      Q => blk00000003_sig00000059
    );
  blk00000003_blk0000000e : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000005c,
      Q => blk00000003_sig0000005d
    );
  blk00000003_blk0000000d : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000005b,
      Q => blk00000003_sig00000057
    );
  blk00000003_blk0000000c : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig0000005a,
      Q => blk00000003_sig00000056
    );
  blk00000003_blk0000000b : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000059,
      Q => blk00000003_sig00000055
    );
  blk00000003_blk0000000a : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000057,
      Q => blk00000003_sig00000058
    );
  blk00000003_blk00000009 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000056,
      Q => blk00000003_sig00000053
    );
  blk00000003_blk00000008 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000055,
      Q => blk00000003_sig00000051
    );
  blk00000003_blk00000007 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000053,
      Q => blk00000003_sig00000054
    );
  blk00000003_blk00000006 : FDE
    generic map(
      INIT => '0'
    )
    port map (
      C => clk,
      CE => ce,
      D => blk00000003_sig00000051,
      Q => blk00000003_sig00000052
    );
  blk00000003_blk00000005 : VCC
    port map (
      P => NlwRenamedSig_OI_rfd
    );
  blk00000003_blk00000004 : GND
    port map (
      G => blk00000003_sig0000004f
    );

end STRUCTURE;

-- synthesis translate_on
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2012 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file mult_11_2_234eb26fa92ee3d2.vhd when simulating
-- the core, mult_11_2_234eb26fa92ee3d2. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY mult_11_2_234eb26fa92ee3d2 IS
  PORT (
    clk : IN STD_LOGIC;
    a : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    ce : IN STD_LOGIC;
    sclr : IN STD_LOGIC;
    p : OUT STD_LOGIC_VECTOR(21 DOWNTO 0)
  );
END mult_11_2_234eb26fa92ee3d2;

ARCHITECTURE mult_11_2_234eb26fa92ee3d2_a OF mult_11_2_234eb26fa92ee3d2 IS
-- synthesis translate_off
COMPONENT wrapped_mult_11_2_234eb26fa92ee3d2
  PORT (
    clk : IN STD_LOGIC;
    a : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    ce : IN STD_LOGIC;
    sclr : IN STD_LOGIC;
    p : OUT STD_LOGIC_VECTOR(21 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_mult_11_2_234eb26fa92ee3d2 USE ENTITY XilinxCoreLib.mult_gen_v11_2(behavioral)
    GENERIC MAP (
      c_a_type => 1,
      c_a_width => 16,
      c_b_type => 1,
      c_b_value => "10000001",
      c_b_width => 6,
      c_ccm_imp => 0,
      c_ce_overrides_sclr => 1,
      c_has_ce => 1,
      c_has_sclr => 1,
      c_has_zero_detect => 0,
      c_latency => 3,
      c_model_type => 0,
      c_mult_type => 1,
      c_optimize_goal => 1,
      c_out_high => 21,
      c_out_low => 0,
      c_round_output => 0,
      c_round_pt => 0,
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_mult_11_2_234eb26fa92ee3d2
  PORT MAP (
    clk => clk,
    a => a,
    b => b,
    ce => ce,
    sclr => sclr,
    p => p
  );
-- synthesis translate_on

END mult_11_2_234eb26fa92ee3d2_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2012 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file mult_11_2_3f458b247f28c718.vhd when simulating
-- the core, mult_11_2_3f458b247f28c718. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY mult_11_2_3f458b247f28c718 IS
  PORT (
    clk : IN STD_LOGIC;
    a : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    ce : IN STD_LOGIC;
    sclr : IN STD_LOGIC;
    p : OUT STD_LOGIC_VECTOR(47 DOWNTO 0)
  );
END mult_11_2_3f458b247f28c718;

ARCHITECTURE mult_11_2_3f458b247f28c718_a OF mult_11_2_3f458b247f28c718 IS
-- synthesis translate_off
COMPONENT wrapped_mult_11_2_3f458b247f28c718
  PORT (
    clk : IN STD_LOGIC;
    a : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    ce : IN STD_LOGIC;
    sclr : IN STD_LOGIC;
    p : OUT STD_LOGIC_VECTOR(47 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_mult_11_2_3f458b247f28c718 USE ENTITY XilinxCoreLib.mult_gen_v11_2(behavioral)
    GENERIC MAP (
      c_a_type => 1,
      c_a_width => 32,
      c_b_type => 1,
      c_b_value => "10000001",
      c_b_width => 16,
      c_ccm_imp => 0,
      c_ce_overrides_sclr => 1,
      c_has_ce => 1,
      c_has_sclr => 1,
      c_has_zero_detect => 0,
      c_latency => 2,
      c_model_type => 0,
      c_mult_type => 1,
      c_optimize_goal => 1,
      c_out_high => 47,
      c_out_low => 0,
      c_round_output => 0,
      c_round_pt => 0,
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_mult_11_2_3f458b247f28c718
  PORT MAP (
    clk => clk,
    a => a,
    b => b,
    ce => ce,
    sclr => sclr,
    p => p
  );
-- synthesis translate_on

END mult_11_2_3f458b247f28c718_a;
--------------------------------------------------------------------------------
--    This file is owned and controlled by Xilinx and must be used solely     --
--    for design, simulation, implementation and creation of design files     --
--    limited to Xilinx devices or technologies. Use with non-Xilinx          --
--    devices or technologies is expressly prohibited and immediately         --
--    terminates your license.                                                --
--                                                                            --
--    XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS" SOLELY    --
--    FOR USE IN DEVELOPING PROGRAMS AND SOLUTIONS FOR XILINX DEVICES.  BY    --
--    PROVIDING THIS DESIGN, CODE, OR INFORMATION AS ONE POSSIBLE             --
--    IMPLEMENTATION OF THIS FEATURE, APPLICATION OR STANDARD, XILINX IS      --
--    MAKING NO REPRESENTATION THAT THIS IMPLEMENTATION IS FREE FROM ANY      --
--    CLAIMS OF INFRINGEMENT, AND YOU ARE RESPONSIBLE FOR OBTAINING ANY       --
--    RIGHTS YOU MAY REQUIRE FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY       --
--    DISCLAIMS ANY WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE   --
--    IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR          --
--    REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF         --
--    INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A   --
--    PARTICULAR PURPOSE.                                                     --
--                                                                            --
--    Xilinx products are not intended for use in life support appliances,    --
--    devices, or systems.  Use in such applications are expressly            --
--    prohibited.                                                             --
--                                                                            --
--    (c) Copyright 1995-2012 Xilinx, Inc.                                    --
--    All rights reserved.                                                    --
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- You must compile the wrapper file mult_11_2_7165ba8b8713bab6.vhd when simulating
-- the core, mult_11_2_7165ba8b8713bab6. When compiling the wrapper file, be sure to
-- reference the XilinxCoreLib VHDL simulation library. For detailed
-- instructions, please refer to the "CORE Generator Help".

-- The synthesis directives "translate_off/translate_on" specified
-- below are supported by Xilinx, Mentor Graphics and Synplicity
-- synthesis tools. Ensure they are correct for your synthesis tool(s).

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
-- synthesis translate_off
LIBRARY XilinxCoreLib;
-- synthesis translate_on
ENTITY mult_11_2_7165ba8b8713bab6 IS
  PORT (
    clk : IN STD_LOGIC;
    a : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    ce : IN STD_LOGIC;
    sclr : IN STD_LOGIC;
    p : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END mult_11_2_7165ba8b8713bab6;

ARCHITECTURE mult_11_2_7165ba8b8713bab6_a OF mult_11_2_7165ba8b8713bab6 IS
-- synthesis translate_off
COMPONENT wrapped_mult_11_2_7165ba8b8713bab6
  PORT (
    clk : IN STD_LOGIC;
    a : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    b : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    ce : IN STD_LOGIC;
    sclr : IN STD_LOGIC;
    p : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
  );
END COMPONENT;

-- Configuration specification
  FOR ALL : wrapped_mult_11_2_7165ba8b8713bab6 USE ENTITY XilinxCoreLib.mult_gen_v11_2(behavioral)
    GENERIC MAP (
      c_a_type => 1,
      c_a_width => 16,
      c_b_type => 1,
      c_b_value => "10000001",
      c_b_width => 16,
      c_ccm_imp => 0,
      c_ce_overrides_sclr => 1,
      c_has_ce => 1,
      c_has_sclr => 1,
      c_has_zero_detect => 0,
      c_latency => 3,
      c_model_type => 0,
      c_mult_type => 1,
      c_optimize_goal => 1,
      c_out_high => 31,
      c_out_low => 0,
      c_round_output => 0,
      c_round_pt => 0,
      c_verbosity => 0,
      c_xdevicefamily => "virtex6"
    );
-- synthesis translate_on
BEGIN
-- synthesis translate_off
U0 : wrapped_mult_11_2_7165ba8b8713bab6
  PORT MAP (
    clk => clk,
    a => a,
    b => b,
    ce => ce,
    sclr => sclr,
    p => p
  );
-- synthesis translate_on

END mult_11_2_7165ba8b8713bab6_a;

-------------------------------------------------------------------
-- System Generator version 13.2 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
package conv_pkg is
    constant simulating : boolean := false
      -- synopsys translate_off
        or true
      -- synopsys translate_on
    ;
    constant xlUnsigned : integer := 1;
    constant xlSigned : integer := 2;
    constant xlWrap : integer := 1;
    constant xlSaturate : integer := 2;
    constant xlTruncate : integer := 1;
    constant xlRound : integer := 2;
    constant xlRoundBanker : integer := 3;
    constant xlAddMode : integer := 1;
    constant xlSubMode : integer := 2;
    attribute black_box : boolean;
    attribute syn_black_box : boolean;
    attribute fpga_dont_touch: string;
    attribute box_type :  string;
    attribute keep : string;
    attribute syn_keep : boolean;
    function std_logic_vector_to_unsigned(inp : std_logic_vector) return unsigned;
    function unsigned_to_std_logic_vector(inp : unsigned) return std_logic_vector;
    function std_logic_vector_to_signed(inp : std_logic_vector) return signed;
    function signed_to_std_logic_vector(inp : signed) return std_logic_vector;
    function unsigned_to_signed(inp : unsigned) return signed;
    function signed_to_unsigned(inp : signed) return unsigned;
    function pos(inp : std_logic_vector; arith : INTEGER) return boolean;
    function all_same(inp: std_logic_vector) return boolean;
    function all_zeros(inp: std_logic_vector) return boolean;
    function is_point_five(inp: std_logic_vector) return boolean;
    function all_ones(inp: std_logic_vector) return boolean;
    function convert_type (inp : std_logic_vector; old_width, old_bin_pt,
                           old_arith, new_width, new_bin_pt, new_arith,
                           quantization, overflow : INTEGER)
        return std_logic_vector;
    function cast (inp : std_logic_vector; old_bin_pt,
                   new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector;
    function vec_slice (inp : std_logic_vector; upper, lower : INTEGER)
        return std_logic_vector;
    function s2u_slice (inp : signed; upper, lower : INTEGER)
        return unsigned;
    function u2u_slice (inp : unsigned; upper, lower : INTEGER)
        return unsigned;
    function s2s_cast (inp : signed; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return signed;
    function u2s_cast (inp : unsigned; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return signed;
    function s2u_cast (inp : signed; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return unsigned;
    function u2u_cast (inp : unsigned; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return unsigned;
    function u2v_cast (inp : unsigned; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return std_logic_vector;
    function s2v_cast (inp : signed; old_bin_pt,
                   new_width, new_bin_pt : INTEGER)
        return std_logic_vector;
    function trunc (inp : std_logic_vector; old_width, old_bin_pt, old_arith,
                    new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector;
    function round_towards_inf (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt,
                                new_arith : INTEGER) return std_logic_vector;
    function round_towards_even (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt,
                                new_arith : INTEGER) return std_logic_vector;
    function max_signed(width : INTEGER) return std_logic_vector;
    function min_signed(width : INTEGER) return std_logic_vector;
    function saturation_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                              old_arith, new_width, new_bin_pt, new_arith
                              : INTEGER) return std_logic_vector;
    function wrap_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                        old_arith, new_width, new_bin_pt, new_arith : INTEGER)
                        return std_logic_vector;
    function fractional_bits(a_bin_pt, b_bin_pt: INTEGER) return INTEGER;
    function integer_bits(a_width, a_bin_pt, b_width, b_bin_pt: INTEGER)
        return INTEGER;
    function sign_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector;
    function zero_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector;
    function zero_ext(inp : std_logic; new_width : INTEGER)
        return std_logic_vector;
    function extend_MSB(inp : std_logic_vector; new_width, arith : INTEGER)
        return std_logic_vector;
    function align_input(inp : std_logic_vector; old_width, delta, new_arith,
                          new_width: INTEGER)
        return std_logic_vector;
    function pad_LSB(inp : std_logic_vector; new_width: integer)
        return std_logic_vector;
    function pad_LSB(inp : std_logic_vector; new_width, arith : integer)
        return std_logic_vector;
    function max(L, R: INTEGER) return INTEGER;
    function min(L, R: INTEGER) return INTEGER;
    function "="(left,right: STRING) return boolean;
    function boolean_to_signed (inp : boolean; width: integer)
        return signed;
    function boolean_to_unsigned (inp : boolean; width: integer)
        return unsigned;
    function boolean_to_vector (inp : boolean)
        return std_logic_vector;
    function std_logic_to_vector (inp : std_logic)
        return std_logic_vector;
    function integer_to_std_logic_vector (inp : integer;  width, arith : integer)
        return std_logic_vector;
    function std_logic_vector_to_integer (inp : std_logic_vector;  arith : integer)
        return integer;
    function std_logic_to_integer(constant inp : std_logic := '0')
        return integer;
    function bin_string_element_to_std_logic_vector (inp : string;  width, index : integer)
        return std_logic_vector;
    function bin_string_to_std_logic_vector (inp : string)
        return std_logic_vector;
    function hex_string_to_std_logic_vector (inp : string; width : integer)
        return std_logic_vector;
    function makeZeroBinStr (width : integer) return STRING;
    function and_reduce(inp: std_logic_vector) return std_logic;
    -- synopsys translate_off
    function is_binary_string_invalid (inp : string)
        return boolean;
    function is_binary_string_undefined (inp : string)
        return boolean;
    function is_XorU(inp : std_logic_vector)
        return boolean;
    function to_real(inp : std_logic_vector; bin_pt : integer; arith : integer)
        return real;
    function std_logic_to_real(inp : std_logic; bin_pt : integer; arith : integer)
        return real;
    function real_to_std_logic_vector (inp : real;  width, bin_pt, arith : integer)
        return std_logic_vector;
    function real_string_to_std_logic_vector (inp : string;  width, bin_pt, arith : integer)
        return std_logic_vector;
    constant display_precision : integer := 20;
    function real_to_string (inp : real) return string;
    function valid_bin_string(inp : string) return boolean;
    function std_logic_vector_to_bin_string(inp : std_logic_vector) return string;
    function std_logic_to_bin_string(inp : std_logic) return string;
    function std_logic_vector_to_bin_string_w_point(inp : std_logic_vector; bin_pt : integer)
        return string;
    function real_to_bin_string(inp : real;  width, bin_pt, arith : integer)
        return string;
    type stdlogic_to_char_t is array(std_logic) of character;
    constant to_char : stdlogic_to_char_t := (
        'U' => 'U',
        'X' => 'X',
        '0' => '0',
        '1' => '1',
        'Z' => 'Z',
        'W' => 'W',
        'L' => 'L',
        'H' => 'H',
        '-' => '-');
    -- synopsys translate_on
end conv_pkg;
package body conv_pkg is
    function std_logic_vector_to_unsigned(inp : std_logic_vector)
        return unsigned
    is
    begin
        return unsigned (inp);
    end;
    function unsigned_to_std_logic_vector(inp : unsigned)
        return std_logic_vector
    is
    begin
        return std_logic_vector(inp);
    end;
    function std_logic_vector_to_signed(inp : std_logic_vector)
        return signed
    is
    begin
        return  signed (inp);
    end;
    function signed_to_std_logic_vector(inp : signed)
        return std_logic_vector
    is
    begin
        return std_logic_vector(inp);
    end;
    function unsigned_to_signed (inp : unsigned)
        return signed
    is
    begin
        return signed(std_logic_vector(inp));
    end;
    function signed_to_unsigned (inp : signed)
        return unsigned
    is
    begin
        return unsigned(std_logic_vector(inp));
    end;
    function pos(inp : std_logic_vector; arith : INTEGER)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        if arith = xlUnsigned then
            return true;
        else
            if vec(width-1) = '0' then
                return true;
            else
                return false;
            end if;
        end if;
        return true;
    end;
    function max_signed(width : INTEGER)
        return std_logic_vector
    is
        variable ones : std_logic_vector(width-2 downto 0);
        variable result : std_logic_vector(width-1 downto 0);
    begin
        ones := (others => '1');
        result(width-1) := '0';
        result(width-2 downto 0) := ones;
        return result;
    end;
    function min_signed(width : INTEGER)
        return std_logic_vector
    is
        variable zeros : std_logic_vector(width-2 downto 0);
        variable result : std_logic_vector(width-1 downto 0);
    begin
        zeros := (others => '0');
        result(width-1) := '1';
        result(width-2 downto 0) := zeros;
        return result;
    end;
    function and_reduce(inp: std_logic_vector) return std_logic
    is
        variable result: std_logic;
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        result := vec(0);
        if width > 1 then
            for i in 1 to width-1 loop
                result := result and vec(i);
            end loop;
        end if;
        return result;
    end;
    function all_same(inp: std_logic_vector) return boolean
    is
        variable result: boolean;
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        result := true;
        if width > 0 then
            for i in 1 to width-1 loop
                if vec(i) /= vec(0) then
                    result := false;
                end if;
            end loop;
        end if;
        return result;
    end;
    function all_zeros(inp: std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable zero : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        zero := (others => '0');
        vec := inp;
        -- synopsys translate_off
        if (is_XorU(vec)) then
            return false;
        end if;
         -- synopsys translate_on
        if (std_logic_vector_to_unsigned(vec) = std_logic_vector_to_unsigned(zero)) then
            result := true;
        else
            result := false;
        end if;
        return result;
    end;
    function is_point_five(inp: std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        vec := inp;
        -- synopsys translate_off
        if (is_XorU(vec)) then
            return false;
        end if;
         -- synopsys translate_on
        if (width > 1) then
           if ((vec(width-1) = '1') and (all_zeros(vec(width-2 downto 0)) = true)) then
               result := true;
           else
               result := false;
           end if;
        else
           if (vec(width-1) = '1') then
               result := true;
           else
               result := false;
           end if;
        end if;
        return result;
    end;
    function all_ones(inp: std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable one : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        one := (others => '1');
        vec := inp;
        -- synopsys translate_off
        if (is_XorU(vec)) then
            return false;
        end if;
         -- synopsys translate_on
        if (std_logic_vector_to_unsigned(vec) = std_logic_vector_to_unsigned(one)) then
            result := true;
        else
            result := false;
        end if;
        return result;
    end;
    function full_precision_num_width(quantization, overflow, old_width,
                                      old_bin_pt, old_arith,
                                      new_width, new_bin_pt, new_arith : INTEGER)
        return integer
    is
        variable result : integer;
    begin
        result := old_width + 2;
        return result;
    end;
    function quantized_num_width(quantization, overflow, old_width, old_bin_pt,
                                 old_arith, new_width, new_bin_pt, new_arith
                                 : INTEGER)
        return integer
    is
        variable right_of_dp, left_of_dp, result : integer;
    begin
        right_of_dp := max(new_bin_pt, old_bin_pt);
        left_of_dp := max((new_width - new_bin_pt), (old_width - old_bin_pt));
        result := (old_width + 2) + (new_bin_pt - old_bin_pt);
        return result;
    end;
    function convert_type (inp : std_logic_vector; old_width, old_bin_pt,
                           old_arith, new_width, new_bin_pt, new_arith,
                           quantization, overflow : INTEGER)
        return std_logic_vector
    is
        constant fp_width : integer :=
            full_precision_num_width(quantization, overflow, old_width,
                                     old_bin_pt, old_arith, new_width,
                                     new_bin_pt, new_arith);
        constant fp_bin_pt : integer := old_bin_pt;
        constant fp_arith : integer := old_arith;
        variable full_precision_result : std_logic_vector(fp_width-1 downto 0);
        constant q_width : integer :=
            quantized_num_width(quantization, overflow, old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt, new_arith);
        constant q_bin_pt : integer := new_bin_pt;
        constant q_arith : integer := old_arith;
        variable quantized_result : std_logic_vector(q_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        result := (others => '0');
        full_precision_result := cast(inp, old_bin_pt, fp_width, fp_bin_pt,
                                      fp_arith);
        if (quantization = xlRound) then
            quantized_result := round_towards_inf(full_precision_result,
                                                  fp_width, fp_bin_pt,
                                                  fp_arith, q_width, q_bin_pt,
                                                  q_arith);
        elsif (quantization = xlRoundBanker) then
            quantized_result := round_towards_even(full_precision_result,
                                                  fp_width, fp_bin_pt,
                                                  fp_arith, q_width, q_bin_pt,
                                                  q_arith);
        else
            quantized_result := trunc(full_precision_result, fp_width, fp_bin_pt,
                                      fp_arith, q_width, q_bin_pt, q_arith);
        end if;
        if (overflow = xlSaturate) then
            result := saturation_arith(quantized_result, q_width, q_bin_pt,
                                       q_arith, new_width, new_bin_pt, new_arith);
        else
             result := wrap_arith(quantized_result, q_width, q_bin_pt, q_arith,
                                  new_width, new_bin_pt, new_arith);
        end if;
        return result;
    end;
    function cast (inp : std_logic_vector; old_bin_pt, new_width,
                   new_bin_pt, new_arith : INTEGER)
        return std_logic_vector
    is
        constant old_width : integer := inp'length;
        constant left_of_dp : integer := (new_width - new_bin_pt)
                                         - (old_width - old_bin_pt);
        constant right_of_dp : integer := (new_bin_pt - old_bin_pt);
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable j   : integer;
    begin
        vec := inp;
        for i in new_width-1 downto 0 loop
            j := i - right_of_dp;
            if ( j > old_width-1) then
                if (new_arith = xlUnsigned) then
                    result(i) := '0';
                else
                    result(i) := vec(old_width-1);
                end if;
            elsif ( j >= 0) then
                result(i) := vec(j);
            else
                result(i) := '0';
            end if;
        end loop;
        return result;
    end;
    function vec_slice (inp : std_logic_vector; upper, lower : INTEGER)
      return std_logic_vector
    is
    begin
        return inp(upper downto lower);
    end;
    function s2u_slice (inp : signed; upper, lower : INTEGER)
      return unsigned
    is
    begin
        return unsigned(vec_slice(std_logic_vector(inp), upper, lower));
    end;
    function u2u_slice (inp : unsigned; upper, lower : INTEGER)
      return unsigned
    is
    begin
        return unsigned(vec_slice(std_logic_vector(inp), upper, lower));
    end;
    function s2s_cast (inp : signed; old_bin_pt, new_width, new_bin_pt : INTEGER)
        return signed
    is
    begin
        return signed(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlSigned));
    end;
    function s2u_cast (inp : signed; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return unsigned
    is
    begin
        return unsigned(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlSigned));
    end;
    function u2s_cast (inp : unsigned; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return signed
    is
    begin
        return signed(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlUnsigned));
    end;
    function u2u_cast (inp : unsigned; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return unsigned
    is
    begin
        return unsigned(cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlUnsigned));
    end;
    function u2v_cast (inp : unsigned; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return std_logic_vector
    is
    begin
        return cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlUnsigned);
    end;
    function s2v_cast (inp : signed; old_bin_pt, new_width,
                   new_bin_pt : INTEGER)
        return std_logic_vector
    is
    begin
        return cast(std_logic_vector(inp), old_bin_pt, new_width, new_bin_pt, xlSigned);
    end;
    function boolean_to_signed (inp : boolean; width : integer)
        return signed
    is
        variable result : signed(width - 1 downto 0);
    begin
        result := (others => '0');
        if inp then
          result(0) := '1';
        else
          result(0) := '0';
        end if;
        return result;
    end;
    function boolean_to_unsigned (inp : boolean; width : integer)
        return unsigned
    is
        variable result : unsigned(width - 1 downto 0);
    begin
        result := (others => '0');
        if inp then
          result(0) := '1';
        else
          result(0) := '0';
        end if;
        return result;
    end;
    function boolean_to_vector (inp : boolean)
        return std_logic_vector
    is
        variable result : std_logic_vector(1 - 1 downto 0);
    begin
        result := (others => '0');
        if inp then
          result(0) := '1';
        else
          result(0) := '0';
        end if;
        return result;
    end;
    function std_logic_to_vector (inp : std_logic)
        return std_logic_vector
    is
        variable result : std_logic_vector(1 - 1 downto 0);
    begin
        result(0) := inp;
        return result;
    end;
    function trunc (inp : std_logic_vector; old_width, old_bin_pt, old_arith,
                                new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector
    is
        constant right_of_dp : integer := (old_bin_pt - new_bin_pt);
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if right_of_dp >= 0 then
            if new_arith = xlUnsigned then
                result := zero_ext(vec(old_width-1 downto right_of_dp), new_width);
            else
                result := sign_ext(vec(old_width-1 downto right_of_dp), new_width);
            end if;
        else
            if new_arith = xlUnsigned then
                result := zero_ext(pad_LSB(vec, old_width +
                                           abs(right_of_dp)), new_width);
            else
                result := sign_ext(pad_LSB(vec, old_width +
                                           abs(right_of_dp)), new_width);
            end if;
        end if;
        return result;
    end;
    function round_towards_inf (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt, new_arith
                                : INTEGER)
        return std_logic_vector
    is
        constant right_of_dp : integer := (old_bin_pt - new_bin_pt);
        constant expected_new_width : integer :=  old_width - right_of_dp  + 1;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable one_or_zero : std_logic_vector(new_width-1 downto 0);
        variable truncated_val : std_logic_vector(new_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if right_of_dp >= 0 then
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            else
                truncated_val := sign_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            end if;
        else
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            else
                truncated_val := sign_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            end if;
        end if;
        one_or_zero := (others => '0');
        if (new_arith = xlSigned) then
            if (vec(old_width-1) = '0') then
                one_or_zero(0) := '1';
            end if;
            if (right_of_dp >= 2) and (right_of_dp <= old_width) then
                if (all_zeros(vec(right_of_dp-2 downto 0)) = false) then
                    one_or_zero(0) := '1';
                end if;
            end if;
            if (right_of_dp >= 1) and (right_of_dp <= old_width) then
                if vec(right_of_dp-1) = '0' then
                    one_or_zero(0) := '0';
                end if;
            else
                one_or_zero(0) := '0';
            end if;
        else
            if (right_of_dp >= 1) and (right_of_dp <= old_width) then
                one_or_zero(0) :=  vec(right_of_dp-1);
            end if;
        end if;
        if new_arith = xlSigned then
            result := signed_to_std_logic_vector(std_logic_vector_to_signed(truncated_val) +
                                                 std_logic_vector_to_signed(one_or_zero));
        else
            result := unsigned_to_std_logic_vector(std_logic_vector_to_unsigned(truncated_val) +
                                                  std_logic_vector_to_unsigned(one_or_zero));
        end if;
        return result;
    end;
    function round_towards_even (inp : std_logic_vector; old_width, old_bin_pt,
                                old_arith, new_width, new_bin_pt, new_arith
                                : INTEGER)
        return std_logic_vector
    is
        constant right_of_dp : integer := (old_bin_pt - new_bin_pt);
        constant expected_new_width : integer :=  old_width - right_of_dp  + 1;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable one_or_zero : std_logic_vector(new_width-1 downto 0);
        variable truncated_val : std_logic_vector(new_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if right_of_dp >= 0 then
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            else
                truncated_val := sign_ext(vec(old_width-1 downto right_of_dp),
                                          new_width);
            end if;
        else
            if new_arith = xlUnsigned then
                truncated_val := zero_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            else
                truncated_val := sign_ext(pad_LSB(vec, old_width +
                                                  abs(right_of_dp)), new_width);
            end if;
        end if;
        one_or_zero := (others => '0');
        if (right_of_dp >= 1) and (right_of_dp <= old_width) then
            if (is_point_five(vec(right_of_dp-1 downto 0)) = false) then
                one_or_zero(0) :=  vec(right_of_dp-1);
            else
                one_or_zero(0) :=  vec(right_of_dp);
            end if;
        end if;
        if new_arith = xlSigned then
            result := signed_to_std_logic_vector(std_logic_vector_to_signed(truncated_val) +
                                                 std_logic_vector_to_signed(one_or_zero));
        else
            result := unsigned_to_std_logic_vector(std_logic_vector_to_unsigned(truncated_val) +
                                                  std_logic_vector_to_unsigned(one_or_zero));
        end if;
        return result;
    end;
    function saturation_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                              old_arith, new_width, new_bin_pt, new_arith
                              : INTEGER)
        return std_logic_vector
    is
        constant left_of_dp : integer := (old_width - old_bin_pt) -
                                         (new_width - new_bin_pt);
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable overflow : boolean;
    begin
        vec := inp;
        overflow := true;
        result := (others => '0');
        if (new_width >= old_width) then
            overflow := false;
        end if;
        if ((old_arith = xlSigned and new_arith = xlSigned) and (old_width > new_width)) then
            if all_same(vec(old_width-1 downto new_width-1)) then
                overflow := false;
            end if;
        end if;
        if (old_arith = xlSigned and new_arith = xlUnsigned) then
            if (old_width > new_width) then
                if all_zeros(vec(old_width-1 downto new_width)) then
                    overflow := false;
                end if;
            else
                if (old_width = new_width) then
                    if (vec(new_width-1) = '0') then
                        overflow := false;
                    end if;
                end if;
            end if;
        end if;
        if (old_arith = xlUnsigned and new_arith = xlUnsigned) then
            if (old_width > new_width) then
                if all_zeros(vec(old_width-1 downto new_width)) then
                    overflow := false;
                end if;
            else
                if (old_width = new_width) then
                    overflow := false;
                end if;
            end if;
        end if;
        if ((old_arith = xlUnsigned and new_arith = xlSigned) and (old_width > new_width)) then
            if all_same(vec(old_width-1 downto new_width-1)) then
                overflow := false;
            end if;
        end if;
        if overflow then
            if new_arith = xlSigned then
                if vec(old_width-1) = '0' then
                    result := max_signed(new_width);
                else
                    result := min_signed(new_width);
                end if;
            else
                if ((old_arith = xlSigned) and vec(old_width-1) = '1') then
                    result := (others => '0');
                else
                    result := (others => '1');
                end if;
            end if;
        else
            if (old_arith = xlSigned) and (new_arith = xlUnsigned) then
                if (vec(old_width-1) = '1') then
                    vec := (others => '0');
                end if;
            end if;
            if new_width <= old_width then
                result := vec(new_width-1 downto 0);
            else
                if new_arith = xlUnsigned then
                    result := zero_ext(vec, new_width);
                else
                    result := sign_ext(vec, new_width);
                end if;
            end if;
        end if;
        return result;
    end;
   function wrap_arith(inp:  std_logic_vector;  old_width, old_bin_pt,
                       old_arith, new_width, new_bin_pt, new_arith : INTEGER)
        return std_logic_vector
    is
        variable result : std_logic_vector(new_width-1 downto 0);
        variable result_arith : integer;
    begin
        if (old_arith = xlSigned) and (new_arith = xlUnsigned) then
            result_arith := xlSigned;
        end if;
        result := cast(inp, old_bin_pt, new_width, new_bin_pt, result_arith);
        return result;
    end;
    function fractional_bits(a_bin_pt, b_bin_pt: INTEGER) return INTEGER is
    begin
        return max(a_bin_pt, b_bin_pt);
    end;
    function integer_bits(a_width, a_bin_pt, b_width, b_bin_pt: INTEGER)
        return INTEGER is
    begin
        return  max(a_width - a_bin_pt, b_width - b_bin_pt);
    end;
    function pad_LSB(inp : std_logic_vector; new_width: integer)
        return STD_LOGIC_VECTOR
    is
        constant orig_width : integer := inp'length;
        variable vec : std_logic_vector(orig_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable pos : integer;
        constant pad_pos : integer := new_width - orig_width - 1;
    begin
        vec := inp;
        pos := new_width-1;
        if (new_width >= orig_width) then
            for i in orig_width-1 downto 0 loop
                result(pos) := vec(i);
                pos := pos - 1;
            end loop;
            if pad_pos >= 0 then
                for i in pad_pos downto 0 loop
                    result(i) := '0';
                end loop;
            end if;
        end if;
        return result;
    end;
    function sign_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector
    is
        constant old_width : integer := inp'length;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if new_width >= old_width then
            result(old_width-1 downto 0) := vec;
            if new_width-1 >= old_width then
                for i in new_width-1 downto old_width loop
                    result(i) := vec(old_width-1);
                end loop;
            end if;
        else
            result(new_width-1 downto 0) := vec(new_width-1 downto 0);
        end if;
        return result;
    end;
    function zero_ext(inp : std_logic_vector; new_width : INTEGER)
        return std_logic_vector
    is
        constant old_width : integer := inp'length;
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if new_width >= old_width then
            result(old_width-1 downto 0) := vec;
            if new_width-1 >= old_width then
                for i in new_width-1 downto old_width loop
                    result(i) := '0';
                end loop;
            end if;
        else
            result(new_width-1 downto 0) := vec(new_width-1 downto 0);
        end if;
        return result;
    end;
    function zero_ext(inp : std_logic; new_width : INTEGER)
        return std_logic_vector
    is
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        result(0) := inp;
        for i in new_width-1 downto 1 loop
            result(i) := '0';
        end loop;
        return result;
    end;
    function extend_MSB(inp : std_logic_vector; new_width, arith : INTEGER)
        return std_logic_vector
    is
        constant orig_width : integer := inp'length;
        variable vec : std_logic_vector(orig_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if arith = xlUnsigned then
            result := zero_ext(vec, new_width);
        else
            result := sign_ext(vec, new_width);
        end if;
        return result;
    end;
    function pad_LSB(inp : std_logic_vector; new_width, arith: integer)
        return STD_LOGIC_VECTOR
    is
        constant orig_width : integer := inp'length;
        variable vec : std_logic_vector(orig_width-1 downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
        variable pos : integer;
    begin
        vec := inp;
        pos := new_width-1;
        if (arith = xlUnsigned) then
            result(pos) := '0';
            pos := pos - 1;
        else
            result(pos) := vec(orig_width-1);
            pos := pos - 1;
        end if;
        if (new_width >= orig_width) then
            for i in orig_width-1 downto 0 loop
                result(pos) := vec(i);
                pos := pos - 1;
            end loop;
            if pos >= 0 then
                for i in pos downto 0 loop
                    result(i) := '0';
                end loop;
            end if;
        end if;
        return result;
    end;
    function align_input(inp : std_logic_vector; old_width, delta, new_arith,
                         new_width: INTEGER)
        return std_logic_vector
    is
        variable vec : std_logic_vector(old_width-1 downto 0);
        variable padded_inp : std_logic_vector((old_width + delta)-1  downto 0);
        variable result : std_logic_vector(new_width-1 downto 0);
    begin
        vec := inp;
        if delta > 0 then
            padded_inp := pad_LSB(vec, old_width+delta);
            result := extend_MSB(padded_inp, new_width, new_arith);
        else
            result := extend_MSB(vec, new_width, new_arith);
        end if;
        return result;
    end;
    function max(L, R: INTEGER) return INTEGER is
    begin
        if L > R then
            return L;
        else
            return R;
        end if;
    end;
    function min(L, R: INTEGER) return INTEGER is
    begin
        if L < R then
            return L;
        else
            return R;
        end if;
    end;
    function "="(left,right: STRING) return boolean is
    begin
        if (left'length /= right'length) then
            return false;
        else
            test : for i in 1 to left'length loop
                if left(i) /= right(i) then
                    return false;
                end if;
            end loop test;
            return true;
        end if;
    end;
    -- synopsys translate_off
    function is_binary_string_invalid (inp : string)
        return boolean
    is
        variable vec : string(1 to inp'length);
        variable result : boolean;
    begin
        vec := inp;
        result := false;
        for i in 1 to vec'length loop
            if ( vec(i) = 'X' ) then
                result := true;
            end if;
        end loop;
        return result;
    end;
    function is_binary_string_undefined (inp : string)
        return boolean
    is
        variable vec : string(1 to inp'length);
        variable result : boolean;
    begin
        vec := inp;
        result := false;
        for i in 1 to vec'length loop
            if ( vec(i) = 'U' ) then
                result := true;
            end if;
        end loop;
        return result;
    end;
    function is_XorU(inp : std_logic_vector)
        return boolean
    is
        constant width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable result : boolean;
    begin
        vec := inp;
        result := false;
        for i in 0 to width-1 loop
            if (vec(i) = 'U') or (vec(i) = 'X') then
                result := true;
            end if;
        end loop;
        return result;
    end;
    function to_real(inp : std_logic_vector; bin_pt : integer; arith : integer)
        return real
    is
        variable  vec : std_logic_vector(inp'length-1 downto 0);
        variable result, shift_val, undefined_real : real;
        variable neg_num : boolean;
    begin
        vec := inp;
        result := 0.0;
        neg_num := false;
        if vec(inp'length-1) = '1' then
            neg_num := true;
        end if;
        for i in 0 to inp'length-1 loop
            if  vec(i) = 'U' or vec(i) = 'X' then
                return undefined_real;
            end if;
            if arith = xlSigned then
                if neg_num then
                    if vec(i) = '0' then
                        result := result + 2.0**i;
                    end if;
                else
                    if vec(i) = '1' then
                        result := result + 2.0**i;
                    end if;
                end if;
            else
                if vec(i) = '1' then
                    result := result + 2.0**i;
                end if;
            end if;
        end loop;
        if arith = xlSigned then
            if neg_num then
                result := result + 1.0;
                result := result * (-1.0);
            end if;
        end if;
        shift_val := 2.0**(-1*bin_pt);
        result := result * shift_val;
        return result;
    end;
    function std_logic_to_real(inp : std_logic; bin_pt : integer; arith : integer)
        return real
    is
        variable result : real := 0.0;
    begin
        if inp = '1' then
            result := 1.0;
        end if;
        if arith = xlSigned then
            assert false
                report "It doesn't make sense to convert a 1 bit number to a signed real.";
        end if;
        return result;
    end;
    -- synopsys translate_on
    function integer_to_std_logic_vector (inp : integer;  width, arith : integer)
        return std_logic_vector
    is
        variable result : std_logic_vector(width-1 downto 0);
        variable unsigned_val : unsigned(width-1 downto 0);
        variable signed_val : signed(width-1 downto 0);
    begin
        if (arith = xlSigned) then
            signed_val := to_signed(inp, width);
            result := signed_to_std_logic_vector(signed_val);
        else
            unsigned_val := to_unsigned(inp, width);
            result := unsigned_to_std_logic_vector(unsigned_val);
        end if;
        return result;
    end;
    function std_logic_vector_to_integer (inp : std_logic_vector;  arith : integer)
        return integer
    is
        constant width : integer := inp'length;
        variable unsigned_val : unsigned(width-1 downto 0);
        variable signed_val : signed(width-1 downto 0);
        variable result : integer;
    begin
        if (arith = xlSigned) then
            signed_val := std_logic_vector_to_signed(inp);
            result := to_integer(signed_val);
        else
            unsigned_val := std_logic_vector_to_unsigned(inp);
            result := to_integer(unsigned_val);
        end if;
        return result;
    end;
    function std_logic_to_integer(constant inp : std_logic := '0')
        return integer
    is
    begin
        if inp = '1' then
            return 1;
        else
            return 0;
        end if;
    end;
    function makeZeroBinStr (width : integer) return STRING is
        variable result : string(1 to width+3);
    begin
        result(1) := '0';
        result(2) := 'b';
        for i in 3 to width+2 loop
            result(i) := '0';
        end loop;
        result(width+3) := '.';
        return result;
    end;
    -- synopsys translate_off
    function real_string_to_std_logic_vector (inp : string;  width, bin_pt, arith : integer)
        return std_logic_vector
    is
        variable result : std_logic_vector(width-1 downto 0);
    begin
        result := (others => '0');
        return result;
    end;
    function real_to_std_logic_vector (inp : real;  width, bin_pt, arith : integer)
        return std_logic_vector
    is
        variable real_val : real;
        variable int_val : integer;
        variable result : std_logic_vector(width-1 downto 0) := (others => '0');
        variable unsigned_val : unsigned(width-1 downto 0) := (others => '0');
        variable signed_val : signed(width-1 downto 0) := (others => '0');
    begin
        real_val := inp;
        int_val := integer(real_val * 2.0**(bin_pt));
        if (arith = xlSigned) then
            signed_val := to_signed(int_val, width);
            result := signed_to_std_logic_vector(signed_val);
        else
            unsigned_val := to_unsigned(int_val, width);
            result := unsigned_to_std_logic_vector(unsigned_val);
        end if;
        return result;
    end;
    -- synopsys translate_on
    function valid_bin_string (inp : string)
        return boolean
    is
        variable vec : string(1 to inp'length);
    begin
        vec := inp;
        if (vec(1) = '0' and vec(2) = 'b') then
            return true;
        else
            return false;
        end if;
    end;
    function hex_string_to_std_logic_vector(inp: string; width : integer)
        return std_logic_vector is
        constant strlen       : integer := inp'LENGTH;
        variable result       : std_logic_vector(width-1 downto 0);
        variable bitval       : std_logic_vector((strlen*4)-1 downto 0);
        variable posn         : integer;
        variable ch           : character;
        variable vec          : string(1 to strlen);
    begin
        vec := inp;
        result := (others => '0');
        posn := (strlen*4)-1;
        for i in 1 to strlen loop
            ch := vec(i);
            case ch is
                when '0' => bitval(posn downto posn-3) := "0000";
                when '1' => bitval(posn downto posn-3) := "0001";
                when '2' => bitval(posn downto posn-3) := "0010";
                when '3' => bitval(posn downto posn-3) := "0011";
                when '4' => bitval(posn downto posn-3) := "0100";
                when '5' => bitval(posn downto posn-3) := "0101";
                when '6' => bitval(posn downto posn-3) := "0110";
                when '7' => bitval(posn downto posn-3) := "0111";
                when '8' => bitval(posn downto posn-3) := "1000";
                when '9' => bitval(posn downto posn-3) := "1001";
                when 'A' | 'a' => bitval(posn downto posn-3) := "1010";
                when 'B' | 'b' => bitval(posn downto posn-3) := "1011";
                when 'C' | 'c' => bitval(posn downto posn-3) := "1100";
                when 'D' | 'd' => bitval(posn downto posn-3) := "1101";
                when 'E' | 'e' => bitval(posn downto posn-3) := "1110";
                when 'F' | 'f' => bitval(posn downto posn-3) := "1111";
                when others => bitval(posn downto posn-3) := "XXXX";
                               -- synopsys translate_off
                               ASSERT false
                                   REPORT "Invalid hex value" SEVERITY ERROR;
                               -- synopsys translate_on
            end case;
            posn := posn - 4;
        end loop;
        if (width <= strlen*4) then
            result :=  bitval(width-1 downto 0);
        else
            result((strlen*4)-1 downto 0) := bitval;
        end if;
        return result;
    end;
    function bin_string_to_std_logic_vector (inp : string)
        return std_logic_vector
    is
        variable pos : integer;
        variable vec : string(1 to inp'length);
        variable result : std_logic_vector(inp'length-1 downto 0);
    begin
        vec := inp;
        pos := inp'length-1;
        result := (others => '0');
        for i in 1 to vec'length loop
            -- synopsys translate_off
            if (pos < 0) and (vec(i) = '0' or vec(i) = '1' or vec(i) = 'X' or vec(i) = 'U')  then
                assert false
                    report "Input string is larger than output std_logic_vector. Truncating output.";
                return result;
            end if;
            -- synopsys translate_on
            if vec(i) = '0' then
                result(pos) := '0';
                pos := pos - 1;
            end if;
            if vec(i) = '1' then
                result(pos) := '1';
                pos := pos - 1;
            end if;
            -- synopsys translate_off
            if (vec(i) = 'X' or vec(i) = 'U') then
                result(pos) := 'U';
                pos := pos - 1;
            end if;
            -- synopsys translate_on
        end loop;
        return result;
    end;
    function bin_string_element_to_std_logic_vector (inp : string;  width, index : integer)
        return std_logic_vector
    is
        constant str_width : integer := width + 4;
        constant inp_len : integer := inp'length;
        constant num_elements : integer := (inp_len + 1)/str_width;
        constant reverse_index : integer := (num_elements-1) - index;
        variable left_pos : integer;
        variable right_pos : integer;
        variable vec : string(1 to inp'length);
        variable result : std_logic_vector(width-1 downto 0);
    begin
        vec := inp;
        result := (others => '0');
        if (reverse_index = 0) and (reverse_index < num_elements) and (inp_len-3 >= width) then
            left_pos := 1;
            right_pos := width + 3;
            result := bin_string_to_std_logic_vector(vec(left_pos to right_pos));
        end if;
        if (reverse_index > 0) and (reverse_index < num_elements) and (inp_len-3 >= width) then
            left_pos := (reverse_index * str_width) + 1;
            right_pos := left_pos + width + 2;
            result := bin_string_to_std_logic_vector(vec(left_pos to right_pos));
        end if;
        return result;
    end;
   -- synopsys translate_off
    function std_logic_vector_to_bin_string(inp : std_logic_vector)
        return string
    is
        variable vec : std_logic_vector(1 to inp'length);
        variable result : string(vec'range);
    begin
        vec := inp;
        for i in vec'range loop
            result(i) := to_char(vec(i));
        end loop;
        return result;
    end;
    function std_logic_to_bin_string(inp : std_logic)
        return string
    is
        variable result : string(1 to 3);
    begin
        result(1) := '0';
        result(2) := 'b';
        result(3) := to_char(inp);
        return result;
    end;
    function std_logic_vector_to_bin_string_w_point(inp : std_logic_vector; bin_pt : integer)
        return string
    is
        variable width : integer := inp'length;
        variable vec : std_logic_vector(width-1 downto 0);
        variable str_pos : integer;
        variable result : string(1 to width+3);
    begin
        vec := inp;
        str_pos := 1;
        result(str_pos) := '0';
        str_pos := 2;
        result(str_pos) := 'b';
        str_pos := 3;
        for i in width-1 downto 0  loop
            if (((width+3) - bin_pt) = str_pos) then
                result(str_pos) := '.';
                str_pos := str_pos + 1;
            end if;
            result(str_pos) := to_char(vec(i));
            str_pos := str_pos + 1;
        end loop;
        if (bin_pt = 0) then
            result(str_pos) := '.';
        end if;
        return result;
    end;
    function real_to_bin_string(inp : real;  width, bin_pt, arith : integer)
        return string
    is
        variable result : string(1 to width);
        variable vec : std_logic_vector(width-1 downto 0);
    begin
        vec := real_to_std_logic_vector(inp, width, bin_pt, arith);
        result := std_logic_vector_to_bin_string(vec);
        return result;
    end;
    function real_to_string (inp : real) return string
    is
        variable result : string(1 to display_precision) := (others => ' ');
    begin
        result(real'image(inp)'range) := real'image(inp);
        return result;
    end;
    -- synopsys translate_on
end conv_pkg;

-------------------------------------------------------------------
-- System Generator version 13.2 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
library thread_id_calc_lib;
use thread_id_calc_lib.conv_pkg.all;
entity srl17e is
    generic (width : integer:=16;
             latency : integer :=8);
    port (clk   : in std_logic;
          ce    : in std_logic;
          d     : in std_logic_vector(width-1 downto 0);
          q     : out std_logic_vector(width-1 downto 0));
end srl17e;
architecture structural of srl17e is
    component SRL16E
        port (D   : in STD_ULOGIC;
              CE  : in STD_ULOGIC;
              CLK : in STD_ULOGIC;
              A0  : in STD_ULOGIC;
              A1  : in STD_ULOGIC;
              A2  : in STD_ULOGIC;
              A3  : in STD_ULOGIC;
              Q   : out STD_ULOGIC);
    end component;
    attribute syn_black_box of SRL16E : component is true;
    attribute fpga_dont_touch of SRL16E : component is "true";
    component FDE
        port(
            Q  :        out   STD_ULOGIC;
            D  :        in    STD_ULOGIC;
            C  :        in    STD_ULOGIC;
            CE :        in    STD_ULOGIC);
    end component;
    attribute syn_black_box of FDE : component is true;
    attribute fpga_dont_touch of FDE : component is "true";
    constant a : std_logic_vector(4 downto 0) :=
        integer_to_std_logic_vector(latency-2,5,xlSigned);
    signal d_delayed : std_logic_vector(width-1 downto 0);
    signal srl16_out : std_logic_vector(width-1 downto 0);
begin
    d_delayed <= d after 200 ps;
    reg_array : for i in 0 to width-1 generate
        srl16_used: if latency > 1 generate
            u1 : srl16e port map(clk => clk,
                                 d => d_delayed(i),
                                 q => srl16_out(i),
                                 ce => ce,
                                 a0 => a(0),
                                 a1 => a(1),
                                 a2 => a(2),
                                 a3 => a(3));
        end generate;
        srl16_not_used: if latency <= 1 generate
            srl16_out(i) <= d_delayed(i);
        end generate;
        fde_used: if latency /= 0  generate
            u2 : fde port map(c => clk,
                              d => srl16_out(i),
                              q => q(i),
                              ce => ce);
        end generate;
        fde_not_used: if latency = 0  generate
            q(i) <= srl16_out(i);
        end generate;
    end generate;
 end structural;
library IEEE;
use IEEE.std_logic_1164.all;
library thread_id_calc_lib;
use thread_id_calc_lib.conv_pkg.all;
entity synth_reg is
    generic (width           : integer := 8;
             latency         : integer := 1);
    port (i       : in std_logic_vector(width-1 downto 0);
          ce      : in std_logic;
          clr     : in std_logic;
          clk     : in std_logic;
          o       : out std_logic_vector(width-1 downto 0));
end synth_reg;
architecture structural of synth_reg is
    component srl17e
        generic (width : integer:=16;
                 latency : integer :=8);
        port (clk : in std_logic;
              ce  : in std_logic;
              d   : in std_logic_vector(width-1 downto 0);
              q   : out std_logic_vector(width-1 downto 0));
    end component;
    function calc_num_srl17es (latency : integer)
        return integer
    is
        variable remaining_latency : integer;
        variable result : integer;
    begin
        result := latency / 17;
        remaining_latency := latency - (result * 17);
        if (remaining_latency /= 0) then
            result := result + 1;
        end if;
        return result;
    end;
    constant complete_num_srl17es : integer := latency / 17;
    constant num_srl17es : integer := calc_num_srl17es(latency);
    constant remaining_latency : integer := latency - (complete_num_srl17es * 17);
    type register_array is array (num_srl17es downto 0) of
        std_logic_vector(width-1 downto 0);
    signal z : register_array;
begin
    z(0) <= i;
    complete_ones : if complete_num_srl17es > 0 generate
        srl17e_array: for i in 0 to complete_num_srl17es-1 generate
            delay_comp : srl17e
                generic map (width => width,
                             latency => 17)
                port map (clk => clk,
                          ce  => ce,
                          d       => z(i),
                          q       => z(i+1));
        end generate;
    end generate;
    partial_one : if remaining_latency > 0 generate
        last_srl17e : srl17e
            generic map (width => width,
                         latency => remaining_latency)
            port map (clk => clk,
                      ce  => ce,
                      d   => z(num_srl17es-1),
                      q   => z(num_srl17es));
    end generate;
    o <= z(num_srl17es);
end structural;
library IEEE;
use IEEE.std_logic_1164.all;
library thread_id_calc_lib;
use thread_id_calc_lib.conv_pkg.all;
entity synth_reg_reg is
    generic (width           : integer := 8;
             latency         : integer := 1);
    port (i       : in std_logic_vector(width-1 downto 0);
          ce      : in std_logic;
          clr     : in std_logic;
          clk     : in std_logic;
          o       : out std_logic_vector(width-1 downto 0));
end synth_reg_reg;
architecture behav of synth_reg_reg is
  type reg_array_type is array (latency-1 downto 0) of std_logic_vector(width -1 downto 0);
  signal reg_bank : reg_array_type := (others => (others => '0'));
  signal reg_bank_in : reg_array_type := (others => (others => '0'));
  attribute syn_allow_retiming : boolean;
  attribute syn_srlstyle : string;
  attribute syn_allow_retiming of reg_bank : signal is true;
  attribute syn_allow_retiming of reg_bank_in : signal is true;
  attribute syn_srlstyle of reg_bank : signal is "registers";
  attribute syn_srlstyle of reg_bank_in : signal is "registers";
begin
  latency_eq_0: if latency = 0 generate
    o <= i;
  end generate latency_eq_0;
  latency_gt_0: if latency >= 1 generate
    o <= reg_bank(latency-1);
    reg_bank_in(0) <= i;
    loop_gen: for idx in latency-2 downto 0 generate
      reg_bank_in(idx+1) <= reg_bank(idx);
    end generate loop_gen;
    sync_loop: for sync_idx in latency-1 downto 0 generate
      sync_proc: process (clk)
      begin
        if clk'event and clk = '1' then
          if ce = '1'  then
            reg_bank(sync_idx) <= reg_bank_in(sync_idx);
          end if;
        end if;
      end process sync_proc;
    end generate sync_loop;
  end generate latency_gt_0;
end behav;

-------------------------------------------------------------------
-- System Generator version 13.2 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
library thread_id_calc_lib;
use thread_id_calc_lib.conv_pkg.all;
entity single_reg_w_init is
  generic (
    width: integer := 8;
    init_index: integer := 0;
    init_value: bit_vector := b"0000"
  );
  port (
    i: in std_logic_vector(width - 1 downto 0);
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    o: out std_logic_vector(width - 1 downto 0)
  );
end single_reg_w_init;
architecture structural of single_reg_w_init is
  function build_init_const(width: integer;
                            init_index: integer;
                            init_value: bit_vector)
    return std_logic_vector
  is
    variable result: std_logic_vector(width - 1 downto 0);
  begin
    if init_index = 0 then
      result := (others => '0');
    elsif init_index = 1 then
      result := (others => '0');
      result(0) := '1';
    else
      result := to_stdlogicvector(init_value);
    end if;
    return result;
  end;
  component fdre
    port (
      q: out std_ulogic;
      d: in  std_ulogic;
      c: in  std_ulogic;
      ce: in  std_ulogic;
      r: in  std_ulogic
    );
  end component;
  attribute syn_black_box of fdre: component is true;
  attribute fpga_dont_touch of fdre: component is "true";
  component fdse
    port (
      q: out std_ulogic;
      d: in  std_ulogic;
      c: in  std_ulogic;
      ce: in  std_ulogic;
      s: in  std_ulogic
    );
  end component;
  attribute syn_black_box of fdse: component is true;
  attribute fpga_dont_touch of fdse: component is "true";
  constant init_const: std_logic_vector(width - 1 downto 0)
    := build_init_const(width, init_index, init_value);
begin
  fd_prim_array: for index in 0 to width - 1 generate
    bit_is_0: if (init_const(index) = '0') generate
      fdre_comp: fdre
        port map (
          c => clk,
          d => i(index),
          q => o(index),
          ce => ce,
          r => clr
        );
    end generate;
    bit_is_1: if (init_const(index) = '1') generate
      fdse_comp: fdse
        port map (
          c => clk,
          d => i(index),
          q => o(index),
          ce => ce,
          s => clr
        );
    end generate;
  end generate;
end architecture structural;
-- synopsys translate_off
library unisim;
use unisim.vcomponents.all;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
library thread_id_calc_lib;
use thread_id_calc_lib.conv_pkg.all;
entity synth_reg_w_init is
  generic (
    width: integer := 8;
    init_index: integer := 0;
    init_value: bit_vector := b"0000";
    latency: integer := 1
  );
  port (
    i: in std_logic_vector(width - 1 downto 0);
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    o: out std_logic_vector(width - 1 downto 0)
  );
end synth_reg_w_init;
architecture structural of synth_reg_w_init is
  component single_reg_w_init
    generic (
      width: integer := 8;
      init_index: integer := 0;
      init_value: bit_vector := b"0000"
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  signal dly_i: std_logic_vector((latency + 1) * width - 1 downto 0);
  signal dly_clr: std_logic;
begin
  latency_eq_0: if (latency = 0) generate
    o <= i;
  end generate;
  latency_gt_0: if (latency >= 1) generate
    dly_i((latency + 1) * width - 1 downto latency * width) <= i
      after 200 ps;
    dly_clr <= clr after 200 ps;
    fd_array: for index in latency downto 1 generate
       reg_comp: single_reg_w_init
          generic map (
            width => width,
            init_index => init_index,
            init_value => init_value
          )
          port map (
            clk => clk,
            i => dly_i((index + 1) * width - 1 downto index * width),
            o => dly_i(index * width - 1 downto (index - 1) * width),
            ce => ce,
            clr => dly_clr
          );
    end generate;
    o <= dly_i(width - 1 downto 0);
  end generate;
end structural;

-------------------------------------------------------------------
-- System Generator version 13.2 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
library thread_id_calc_lib;
use thread_id_calc_lib.conv_pkg.all;
entity xladdsub is
  generic (
    core_name0: string := "";
    a_width: integer := 16;
    a_bin_pt: integer := 4;
    a_arith: integer := xlUnsigned;
    c_in_width: integer := 16;
    c_in_bin_pt: integer := 4;
    c_in_arith: integer := xlUnsigned;
    c_out_width: integer := 16;
    c_out_bin_pt: integer := 4;
    c_out_arith: integer := xlUnsigned;
    b_width: integer := 8;
    b_bin_pt: integer := 2;
    b_arith: integer := xlUnsigned;
    s_width: integer := 17;
    s_bin_pt: integer := 4;
    s_arith: integer := xlUnsigned;
    rst_width: integer := 1;
    rst_bin_pt: integer := 0;
    rst_arith: integer := xlUnsigned;
    en_width: integer := 1;
    en_bin_pt: integer := 0;
    en_arith: integer := xlUnsigned;
    full_s_width: integer := 17;
    full_s_arith: integer := xlUnsigned;
    mode: integer := xlAddMode;
    extra_registers: integer := 0;
    latency: integer := 0;
    quantization: integer := xlTruncate;
    overflow: integer := xlWrap;
    c_latency: integer := 0;
    c_output_width: integer := 17;
    c_has_c_in : integer := 0;
    c_has_c_out : integer := 0
  );
  port (
    a: in std_logic_vector(a_width - 1 downto 0);
    b: in std_logic_vector(b_width - 1 downto 0);
    c_in : in std_logic_vector (0 downto 0) := "0";
    ce: in std_logic;
    clr: in std_logic := '0';
    clk: in std_logic;
    rst: in std_logic_vector(rst_width - 1 downto 0) := "0";
    en: in std_logic_vector(en_width - 1 downto 0) := "1";
    c_out : out std_logic_vector (0 downto 0);
    s: out std_logic_vector(s_width - 1 downto 0)
  );
end xladdsub;
architecture behavior of xladdsub is
  component synth_reg
    generic (
      width: integer := 16;
      latency: integer := 5
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  function format_input(inp: std_logic_vector; old_width, delta, new_arith,
                        new_width: integer)
    return std_logic_vector
  is
    variable vec: std_logic_vector(old_width-1 downto 0);
    variable padded_inp: std_logic_vector((old_width + delta)-1  downto 0);
    variable result: std_logic_vector(new_width-1 downto 0);
  begin
    vec := inp;
    if (delta > 0) then
      padded_inp := pad_LSB(vec, old_width+delta);
      result := extend_MSB(padded_inp, new_width, new_arith);
    else
      result := extend_MSB(vec, new_width, new_arith);
    end if;
    return result;
  end;
  constant full_s_bin_pt: integer := fractional_bits(a_bin_pt, b_bin_pt);
  constant full_a_width: integer := full_s_width;
  constant full_b_width: integer := full_s_width;
  signal full_a: std_logic_vector(full_a_width - 1 downto 0);
  signal full_b: std_logic_vector(full_b_width - 1 downto 0);
  signal core_s: std_logic_vector(full_s_width - 1 downto 0);
  signal conv_s: std_logic_vector(s_width - 1 downto 0);
  signal temp_cout : std_logic;
  signal internal_clr: std_logic;
  signal internal_ce: std_logic;
  signal extra_reg_ce: std_logic;
  signal override: std_logic;
  signal logic1: std_logic_vector(0 downto 0);
  component addsb_11_0_f45daeb7eb283db0
    port (
          a: in std_logic_vector(33 - 1 downto 0);
    s: out std_logic_vector(c_output_width - 1 downto 0);
    b: in std_logic_vector(33 - 1 downto 0)
    );
  end component;
  attribute syn_black_box of addsb_11_0_f45daeb7eb283db0:
    component is true;
  attribute fpga_dont_touch of addsb_11_0_f45daeb7eb283db0:
    component is "true";
  attribute box_type of addsb_11_0_f45daeb7eb283db0:
    component  is "black_box";
begin
  internal_clr <= (clr or (rst(0))) and ce;
  internal_ce <= ce and en(0);
  logic1(0) <= '1';
  addsub_process: process (a, b, core_s)
  begin
    full_a <= format_input (a, a_width, b_bin_pt - a_bin_pt, a_arith,
                            full_a_width);
    full_b <= format_input (b, b_width, a_bin_pt - b_bin_pt, b_arith,
                            full_b_width);
    conv_s <= convert_type (core_s, full_s_width, full_s_bin_pt, full_s_arith,
                            s_width, s_bin_pt, s_arith, quantization, overflow);
  end process addsub_process;

  comp0: if ((core_name0 = "addsb_11_0_f45daeb7eb283db0")) generate
    core_instance0: addsb_11_0_f45daeb7eb283db0
      port map (
         a => full_a,
         s => core_s,
         b => full_b
      );
  end generate;
  latency_test: if (extra_registers > 0) generate
      override_test: if (c_latency > 1) generate
       override_pipe: synth_reg
          generic map (
            width => 1,
            latency => c_latency
          )
          port map (
            i => logic1,
            ce => internal_ce,
            clr => internal_clr,
            clk => clk,
            o(0) => override);
       extra_reg_ce <= ce and en(0) and override;
      end generate override_test;
      no_override: if ((c_latency = 0) or (c_latency = 1)) generate
       extra_reg_ce <= ce and en(0);
      end generate no_override;
      extra_reg: synth_reg
        generic map (
          width => s_width,
          latency => extra_registers
        )
        port map (
          i => conv_s,
          ce => extra_reg_ce,
          clr => internal_clr,
          clk => clk,
          o => s
        );
      cout_test: if (c_has_c_out = 1) generate
      c_out_extra_reg: synth_reg
        generic map (
          width => 1,
          latency => extra_registers
        )
        port map (
          i(0) => temp_cout,
          ce => extra_reg_ce,
          clr => internal_clr,
          clk => clk,
          o => c_out
        );
      end generate cout_test;
  end generate;
  latency_s: if ((latency = 0) or (extra_registers = 0)) generate
    s <= conv_s;
  end generate latency_s;
  latency0: if (((latency = 0) or (extra_registers = 0)) and
                 (c_has_c_out = 1)) generate
    c_out(0) <= temp_cout;
  end generate latency0;
  tie_dangling_cout: if (c_has_c_out = 0) generate
    c_out <= "0";
  end generate tie_dangling_cout;
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library thread_id_calc_lib;
use thread_id_calc_lib.conv_pkg.all;

entity constant_7db069ad14 is
  port (
    op : out std_logic_vector((8 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end constant_7db069ad14;


architecture behavior of constant_7db069ad14 is
begin
  op <= "00110000";
end behavior;


-------------------------------------------------------------------
-- System Generator version 13.2 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
library thread_id_calc_lib;
use thread_id_calc_lib.conv_pkg.all;
entity convert_func_call is
    generic (
        din_width    : integer := 16;
        din_bin_pt   : integer := 4;
        din_arith    : integer := xlUnsigned;
        dout_width   : integer := 8;
        dout_bin_pt  : integer := 2;
        dout_arith   : integer := xlUnsigned;
        quantization : integer := xlTruncate;
        overflow     : integer := xlWrap);
    port (
        din : in std_logic_vector (din_width-1 downto 0);
        result : out std_logic_vector (dout_width-1 downto 0));
end convert_func_call;
architecture behavior of convert_func_call is
begin
    result <= convert_type(din, din_width, din_bin_pt, din_arith,
                           dout_width, dout_bin_pt, dout_arith,
                           quantization, overflow);
end behavior;
library IEEE;
use IEEE.std_logic_1164.all;
library thread_id_calc_lib;
use thread_id_calc_lib.conv_pkg.all;
entity xlconvert is
    generic (
        din_width    : integer := 16;
        din_bin_pt   : integer := 4;
        din_arith    : integer := xlUnsigned;
        dout_width   : integer := 8;
        dout_bin_pt  : integer := 2;
        dout_arith   : integer := xlUnsigned;
        en_width     : integer := 1;
        en_bin_pt    : integer := 0;
        en_arith     : integer := xlUnsigned;
        bool_conversion : integer :=0;
        latency      : integer := 0;
        quantization : integer := xlTruncate;
        overflow     : integer := xlWrap);
    port (
        din : in std_logic_vector (din_width-1 downto 0);
        en  : in std_logic_vector (en_width-1 downto 0);
        ce  : in std_logic;
        clr : in std_logic;
        clk : in std_logic;
        dout : out std_logic_vector (dout_width-1 downto 0));
end xlconvert;
architecture behavior of xlconvert is
    component synth_reg
        generic (width       : integer;
                 latency     : integer);
        port (i       : in std_logic_vector(width-1 downto 0);
              ce      : in std_logic;
              clr     : in std_logic;
              clk     : in std_logic;
              o       : out std_logic_vector(width-1 downto 0));
    end component;
    component convert_func_call
        generic (
            din_width    : integer := 16;
            din_bin_pt   : integer := 4;
            din_arith    : integer := xlUnsigned;
            dout_width   : integer := 8;
            dout_bin_pt  : integer := 2;
            dout_arith   : integer := xlUnsigned;
            quantization : integer := xlTruncate;
            overflow     : integer := xlWrap);
        port (
            din : in std_logic_vector (din_width-1 downto 0);
            result : out std_logic_vector (dout_width-1 downto 0));
    end component;
    -- synopsys translate_off
    -- synopsys translate_on
    signal result : std_logic_vector(dout_width-1 downto 0);
    signal internal_ce : std_logic;
begin
    -- synopsys translate_off
    -- synopsys translate_on
    internal_ce <= ce and en(0);

    bool_conversion_generate : if (bool_conversion = 1)
    generate
      result <= din;
    end generate;
    std_conversion_generate : if (bool_conversion = 0)
    generate
      convert : convert_func_call
        generic map (
          din_width   => din_width,
          din_bin_pt  => din_bin_pt,
          din_arith   => din_arith,
          dout_width  => dout_width,
          dout_bin_pt => dout_bin_pt,
          dout_arith  => dout_arith,
          quantization => quantization,
          overflow     => overflow)
        port map (
          din => din,
          result => result);
    end generate;
    latency_test : if (latency > 0) generate
        reg : synth_reg
            generic map (
              width => dout_width,
              latency => latency
            )
            port map (
              i => result,
              ce => internal_ce,
              clr => clr,
              clk => clk,
              o => dout
            );
    end generate;
    latency0 : if (latency = 0)
    generate
        dout <= result;
    end generate latency0;
end  behavior;

-------------------------------------------------------------------
-- System Generator version 13.2 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
library thread_id_calc_lib;
use thread_id_calc_lib.conv_pkg.all;
entity xlcounter_free is
  generic (
    core_name0: string := "";
    op_width: integer := 5;
    op_arith: integer := xlSigned
  );
  port (
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    op: out std_logic_vector(op_width - 1 downto 0);
    up: in std_logic_vector(0 downto 0) := (others => '0');
    load: in std_logic_vector(0 downto 0) := (others => '0');
    din: in std_logic_vector(op_width - 1 downto 0) := (others => '0');
    en: in std_logic_vector(0 downto 0);
    rst: in std_logic_vector(0 downto 0)
  );
end xlcounter_free ;
architecture behavior of xlcounter_free is
  component cntr_11_0_e7514e290b172ea1
    port (
      clk: in std_logic;
      ce: in std_logic;
      SINIT: in std_logic;
      q: out std_logic_vector(op_width - 1 downto 0)
    );
  end component;
  attribute syn_black_box of cntr_11_0_e7514e290b172ea1:
    component is true;
  attribute fpga_dont_touch of cntr_11_0_e7514e290b172ea1:
    component is "true";
  attribute box_type of cntr_11_0_e7514e290b172ea1:
    component  is "black_box";
-- synopsys translate_off
  constant zeroVec: std_logic_vector(op_width - 1 downto 0) := (others => '0');
  constant oneVec: std_logic_vector(op_width - 1 downto 0) := (others => '1');
  constant zeroStr: string(1 to op_width) :=
    std_logic_vector_to_bin_string(zeroVec);
  constant oneStr: string(1 to op_width) :=
    std_logic_vector_to_bin_string(oneVec);
-- synopsys translate_on
  signal core_sinit: std_logic;
  signal core_ce: std_logic;
  signal op_net: std_logic_vector(op_width - 1 downto 0);
begin
  core_ce <= ce and en(0);
  core_sinit <= (clr or rst(0)) and ce;
  op <= op_net;
  comp0: if ((core_name0 = "cntr_11_0_e7514e290b172ea1")) generate
    core_instance0: cntr_11_0_e7514e290b172ea1
      port map (
        clk => clk,
        ce => core_ce,
        SINIT => core_sinit,
        q => op_net
      );
  end generate;
end behavior;

-------------------------------------------------------------------
-- System Generator version 13.2 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
library thread_id_calc_lib;
use thread_id_calc_lib.conv_pkg.all;
entity xldelay is
   generic(width        : integer := -1;
           latency      : integer := -1;
           reg_retiming : integer := 0);
   port(d       : in std_logic_vector (width-1 downto 0);
        ce      : in std_logic;
        clk     : in std_logic;
        en      : in std_logic;
        q       : out std_logic_vector (width-1 downto 0));
end xldelay;
architecture behavior of xldelay is
   component synth_reg
      generic (width       : integer;
               latency     : integer);
      port (i       : in std_logic_vector(width-1 downto 0);
            ce      : in std_logic;
            clr     : in std_logic;
            clk     : in std_logic;
            o       : out std_logic_vector(width-1 downto 0));
   end component;
   component synth_reg_reg
      generic (width       : integer;
               latency     : integer);
      port (i       : in std_logic_vector(width-1 downto 0);
            ce      : in std_logic;
            clr     : in std_logic;
            clk     : in std_logic;
            o       : out std_logic_vector(width-1 downto 0));
   end component;
   signal internal_ce  : std_logic;
begin
   internal_ce  <= ce and en;
   srl_delay: if (reg_retiming = 0) or (latency < 1) generate
     synth_reg_srl_inst : synth_reg
       generic map (
         width   => width,
         latency => latency)
       port map (
         i   => d,
         ce  => internal_ce,
         clr => '0',
         clk => clk,
         o   => q);
   end generate srl_delay;
   reg_delay: if (reg_retiming = 1) and (latency >= 1) generate
     synth_reg_reg_inst : synth_reg_reg
       generic map (
         width   => width,
         latency => latency)
       port map (
         i   => d,
         ce  => internal_ce,
         clr => '0',
         clk => clk,
         o   => q);
   end generate reg_delay;
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library thread_id_calc_lib;
use thread_id_calc_lib.conv_pkg.all;

entity logical_0d8e48dd8a is
  port (
    d0 : in std_logic_vector((16 - 1) downto 0);
    d1 : in std_logic_vector((32 - 1) downto 0);
    d2 : in std_logic_vector((32 - 1) downto 0);
    y : out std_logic_vector((32 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end logical_0d8e48dd8a;


architecture behavior of logical_0d8e48dd8a is
  signal d0_1_24: std_logic_vector((16 - 1) downto 0);
  signal d1_1_27: std_logic_vector((32 - 1) downto 0);
  signal d2_1_30: std_logic_vector((32 - 1) downto 0);
  signal cast_convert_2_19: std_logic_vector((32 - 1) downto 0);
  signal fully_2_1_bit: std_logic_vector((32 - 1) downto 0);
begin
  d0_1_24 <= d0;
  d1_1_27 <= d1;
  d2_1_30 <= d2;
  cast_convert_2_19 <= cast(d0_1_24, 0, 32, 0, xlUnsigned);
  fully_2_1_bit <= cast_convert_2_19 or d1_1_27 or d2_1_30;
  y <= fully_2_1_bit;
end behavior;


-------------------------------------------------------------------
-- System Generator version 13.2 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
-- synopsys translate_off
library XilinxCoreLib;
-- synopsys translate_on
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
library thread_id_calc_lib;
use thread_id_calc_lib.conv_pkg.all;
entity xlmult is
  generic (
    core_name0: string := "";
    a_width: integer := 4;
    a_bin_pt: integer := 2;
    a_arith: integer := xlSigned;
    b_width: integer := 4;
    b_bin_pt: integer := 1;
    b_arith: integer := xlSigned;
    p_width: integer := 8;
    p_bin_pt: integer := 2;
    p_arith: integer := xlSigned;
    rst_width: integer := 1;
    rst_bin_pt: integer := 0;
    rst_arith: integer := xlUnsigned;
    en_width: integer := 1;
    en_bin_pt: integer := 0;
    en_arith: integer := xlUnsigned;
    quantization: integer := xlTruncate;
    overflow: integer := xlWrap;
    extra_registers: integer := 0;
    c_a_width: integer := 7;
    c_b_width: integer := 7;
    c_type: integer := 0;
    c_a_type: integer := 0;
    c_b_type: integer := 0;
    c_pipelined: integer := 1;
    c_baat: integer := 4;
    multsign: integer := xlSigned;
    c_output_width: integer := 16
  );
  port (
    a: in std_logic_vector(a_width - 1 downto 0);
    b: in std_logic_vector(b_width - 1 downto 0);
    ce: in std_logic;
    clr: in std_logic;
    clk: in std_logic;
    core_ce: in std_logic := '0';
    core_clr: in std_logic := '0';
    core_clk: in std_logic := '0';
    rst: in std_logic_vector(rst_width - 1 downto 0);
    en: in std_logic_vector(en_width - 1 downto 0);
    p: out std_logic_vector(p_width - 1 downto 0)
  );
end xlmult;
architecture behavior of xlmult is
  component synth_reg
    generic (
      width: integer := 16;
      latency: integer := 5
    );
    port (
      i: in std_logic_vector(width - 1 downto 0);
      ce: in std_logic;
      clr: in std_logic;
      clk: in std_logic;
      o: out std_logic_vector(width - 1 downto 0)
    );
  end component;
  component mult_11_2_7165ba8b8713bab6
    port (
      b: in std_logic_vector(c_b_width - 1 downto 0);
      p: out std_logic_vector(c_output_width - 1 downto 0);
      clk: in std_logic;
      ce: in std_logic;
      sclr: in std_logic;
      a: in std_logic_vector(c_a_width - 1 downto 0)
    );
  end component;
  attribute syn_black_box of mult_11_2_7165ba8b8713bab6:
    component is true;
  attribute fpga_dont_touch of mult_11_2_7165ba8b8713bab6:
    component is "true";
  attribute box_type of mult_11_2_7165ba8b8713bab6:
    component  is "black_box";
  component mult_11_2_3f458b247f28c718
    port (
      b: in std_logic_vector(c_b_width - 1 downto 0);
      p: out std_logic_vector(c_output_width - 1 downto 0);
      clk: in std_logic;
      ce: in std_logic;
      sclr: in std_logic;
      a: in std_logic_vector(c_a_width - 1 downto 0)
    );
  end component;
  attribute syn_black_box of mult_11_2_3f458b247f28c718:
    component is true;
  attribute fpga_dont_touch of mult_11_2_3f458b247f28c718:
    component is "true";
  attribute box_type of mult_11_2_3f458b247f28c718:
    component  is "black_box";
  component mult_11_2_234eb26fa92ee3d2
    port (
      b: in std_logic_vector(c_b_width - 1 downto 0);
      p: out std_logic_vector(c_output_width - 1 downto 0);
      clk: in std_logic;
      ce: in std_logic;
      sclr: in std_logic;
      a: in std_logic_vector(c_a_width - 1 downto 0)
    );
  end component;
  attribute syn_black_box of mult_11_2_234eb26fa92ee3d2:
    component is true;
  attribute fpga_dont_touch of mult_11_2_234eb26fa92ee3d2:
    component is "true";
  attribute box_type of mult_11_2_234eb26fa92ee3d2:
    component  is "black_box";
  signal tmp_a: std_logic_vector(c_a_width - 1 downto 0);
  signal conv_a: std_logic_vector(c_a_width - 1 downto 0);
  signal tmp_b: std_logic_vector(c_b_width - 1 downto 0);
  signal conv_b: std_logic_vector(c_b_width - 1 downto 0);
  signal tmp_p: std_logic_vector(c_output_width - 1 downto 0);
  signal conv_p: std_logic_vector(p_width - 1 downto 0);
  -- synopsys translate_off
  signal real_a, real_b, real_p: real;
  -- synopsys translate_on
  signal rfd: std_logic;
  signal rdy: std_logic;
  signal nd: std_logic;
  signal internal_ce: std_logic;
  signal internal_clr: std_logic;
  signal internal_core_ce: std_logic;
begin
-- synopsys translate_off
-- synopsys translate_on
  internal_ce <= ce and en(0);
  internal_core_ce <= core_ce and en(0);
  internal_clr <= (clr or rst(0)) and ce;
  nd <= internal_ce;
  input_process:  process (a,b)
  begin
    tmp_a <= zero_ext(a, c_a_width);
    tmp_b <= zero_ext(b, c_b_width);
  end process;
  output_process: process (tmp_p)
  begin
    conv_p <= convert_type(tmp_p, c_output_width, a_bin_pt+b_bin_pt, multsign,
                           p_width, p_bin_pt, p_arith, quantization, overflow);
  end process;
  comp0: if ((core_name0 = "mult_11_2_7165ba8b8713bab6")) generate
    core_instance0: mult_11_2_7165ba8b8713bab6
      port map (
        a => tmp_a,
        clk => clk,
        ce => internal_ce,
        sclr => internal_clr,
        p => tmp_p,
        b => tmp_b
      );
  end generate;
  comp1: if ((core_name0 = "mult_11_2_3f458b247f28c718")) generate
    core_instance1: mult_11_2_3f458b247f28c718
      port map (
        a => tmp_a,
        clk => clk,
        ce => internal_ce,
        sclr => internal_clr,
        p => tmp_p,
        b => tmp_b
      );
  end generate;
  comp2: if ((core_name0 = "mult_11_2_234eb26fa92ee3d2")) generate
    core_instance2: mult_11_2_234eb26fa92ee3d2
      port map (
        a => tmp_a,
        clk => clk,
        ce => internal_ce,
        sclr => internal_clr,
        p => tmp_p,
        b => tmp_b
      );
  end generate;
  latency_gt_0: if (extra_registers > 0) generate
    reg: synth_reg
      generic map (
        width => p_width,
        latency => extra_registers
      )
      port map (
        i => conv_p,
        ce => internal_ce,
        clr => internal_clr,
        clk => clk,
        o => p
      );
  end generate;
  latency_eq_0: if (extra_registers = 0) generate
    p <= conv_p;
  end generate;
end architecture behavior;

-------------------------------------------------------------------
-- System Generator version 13.2 VHDL source file.
--
-- Copyright(C) 2011 by Xilinx, Inc.  All rights reserved.  This
-- text/file contains proprietary, confidential information of Xilinx,
-- Inc., is distributed under license from Xilinx, Inc., and may be used,
-- copied and/or disclosed only pursuant to the terms of a valid license
-- agreement with Xilinx, Inc.  Xilinx hereby grants you a license to use
-- this text/file solely for design, simulation, implementation and
-- creation of design files limited to Xilinx devices or technologies.
-- Use with non-Xilinx devices or technologies is expressly prohibited
-- and immediately terminates your license unless covered by a separate
-- agreement.
--
-- Xilinx is providing this design, code, or information "as is" solely
-- for use in developing programs and solutions for Xilinx devices.  By
-- providing this design, code, or information as one possible
-- implementation of this feature, application or standard, Xilinx is
-- making no representation that this implementation is free from any
-- claims of infringement.  You are responsible for obtaining any rights
-- you may require for your implementation.  Xilinx expressly disclaims
-- any warranty whatsoever with respect to the adequacy of the
-- implementation, including but not limited to warranties of
-- merchantability or fitness for a particular purpose.
--
-- Xilinx products are not intended for use in life support appliances,
-- devices, or systems.  Use in such applications is expressly prohibited.
--
-- Any modifications that are made to the source code are done at the user's
-- sole risk and will be unsupported.
--
-- This copyright and support notice must be retained as part of this
-- text at all times.  (c) Copyright 1995-2011 Xilinx, Inc.  All rights
-- reserved.
-------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
library thread_id_calc_lib;
use thread_id_calc_lib.conv_pkg.all;
entity xlregister is
   generic (d_width          : integer := 5;
            init_value       : bit_vector := b"00");
   port (d   : in std_logic_vector (d_width-1 downto 0);
         rst : in std_logic_vector(0 downto 0) := "0";
         en  : in std_logic_vector(0 downto 0) := "1";
         ce  : in std_logic;
         clk : in std_logic;
         q   : out std_logic_vector (d_width-1 downto 0));
end xlregister;
architecture behavior of xlregister is
   component synth_reg_w_init
      generic (width      : integer;
               init_index : integer;
               init_value : bit_vector;
               latency    : integer);
      port (i   : in std_logic_vector(width-1 downto 0);
            ce  : in std_logic;
            clr : in std_logic;
            clk : in std_logic;
            o   : out std_logic_vector(width-1 downto 0));
   end component;
   -- synopsys translate_off
   signal real_d, real_q           : real;
   -- synopsys translate_on
   signal internal_clr             : std_logic;
   signal internal_ce              : std_logic;
begin
   internal_clr <= rst(0) and ce;
   internal_ce  <= en(0) and ce;
   synth_reg_inst : synth_reg_w_init
      generic map (width      => d_width,
                   init_index => 2,
                   init_value => init_value,
                   latency    => 1)
      port map (i   => d,
                ce  => internal_ce,
                clr => internal_clr,
                clk => clk,
                o   => q);
end architecture behavior;
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library thread_id_calc_lib;
use thread_id_calc_lib.conv_pkg.all;

entity relational_54048c8b02 is
  port (
    a : in std_logic_vector((8 - 1) downto 0);
    b : in std_logic_vector((8 - 1) downto 0);
    op : out std_logic_vector((1 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end relational_54048c8b02;


architecture behavior of relational_54048c8b02 is
  signal a_1_31: unsigned((8 - 1) downto 0);
  signal b_1_34: unsigned((8 - 1) downto 0);
  signal result_12_3_rel: boolean;
begin
  a_1_31 <= std_logic_vector_to_unsigned(a);
  b_1_34 <= std_logic_vector_to_unsigned(b);
  result_12_3_rel <= a_1_31 = b_1_34;
  op <= boolean_to_vector(result_12_3_rel);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library thread_id_calc_lib;
use thread_id_calc_lib.conv_pkg.all;

entity shift_63b52ec892 is
  port (
    ip : in std_logic_vector((16 - 1) downto 0);
    op : out std_logic_vector((32 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end shift_63b52ec892;


architecture behavior of shift_63b52ec892 is
  signal ip_1_23: unsigned((16 - 1) downto 0);
  type array_type_op_mem_46_20 is array (0 to (1 - 1)) of unsigned((32 - 1) downto 0);
  signal op_mem_46_20: array_type_op_mem_46_20 := (
    0 => "00000000000000000000000000000000");
  signal op_mem_46_20_front_din: unsigned((32 - 1) downto 0);
  signal op_mem_46_20_back: unsigned((32 - 1) downto 0);
  signal op_mem_46_20_push_front_pop_back_en: std_logic;
  signal cast_internal_ip_25_3_lsh: unsigned((42 - 1) downto 0);
  signal internal_ip_33_3_convert: unsigned((32 - 1) downto 0);
begin
  ip_1_23 <= std_logic_vector_to_unsigned(ip);
  op_mem_46_20_back <= op_mem_46_20(0);
  proc_op_mem_46_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_46_20_push_front_pop_back_en = '1')) then
        op_mem_46_20(0) <= op_mem_46_20_front_din;
      end if;
    end if;
  end process proc_op_mem_46_20;
  cast_internal_ip_25_3_lsh <= u2u_cast(ip_1_23, 0, 42, 26);
  internal_ip_33_3_convert <= std_logic_vector_to_unsigned(convert_type(unsigned_to_std_logic_vector(cast_internal_ip_25_3_lsh), 42, 0, xlUnsigned, 32, 0, xlUnsigned, xlTruncate, xlSaturate));
  op_mem_46_20_push_front_pop_back_en <= '0';
  op <= unsigned_to_std_logic_vector(internal_ip_33_3_convert);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library thread_id_calc_lib;
use thread_id_calc_lib.conv_pkg.all;

entity shift_cdf6c3fa1e is
  port (
    ip : in std_logic_vector((16 - 1) downto 0);
    op : out std_logic_vector((32 - 1) downto 0);
    clk : in std_logic;
    ce : in std_logic;
    clr : in std_logic);
end shift_cdf6c3fa1e;


architecture behavior of shift_cdf6c3fa1e is
  signal ip_1_23: unsigned((16 - 1) downto 0);
  type array_type_op_mem_46_20 is array (0 to (1 - 1)) of unsigned((32 - 1) downto 0);
  signal op_mem_46_20: array_type_op_mem_46_20 := (
    0 => "00000000000000000000000000000000");
  signal op_mem_46_20_front_din: unsigned((32 - 1) downto 0);
  signal op_mem_46_20_back: unsigned((32 - 1) downto 0);
  signal op_mem_46_20_push_front_pop_back_en: std_logic;
  signal cast_internal_ip_25_3_lsh: unsigned((32 - 1) downto 0);
begin
  ip_1_23 <= std_logic_vector_to_unsigned(ip);
  op_mem_46_20_back <= op_mem_46_20(0);
  proc_op_mem_46_20: process (clk)
  is
    variable i: integer;
  begin
    if (clk'event and (clk = '1')) then
      if ((ce = '1') and (op_mem_46_20_push_front_pop_back_en = '1')) then
        op_mem_46_20(0) <= op_mem_46_20_front_din;
      end if;
    end if;
  end process proc_op_mem_46_20;
  cast_internal_ip_25_3_lsh <= u2u_cast(ip_1_23, 0, 32, 16);
  op_mem_46_20_push_front_pop_back_en <= '0';
  op <= unsigned_to_std_logic_vector(cast_internal_ip_25_3_lsh);
end behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library thread_id_calc_lib;
use thread_id_calc_lib.conv_pkg.all;

entity xldivider_generator_4c82698e6ec63d36ca8d57faf12d4ed2 is 
  port(
    ce:in std_logic;
    clk:in std_logic;
    dividend:in std_logic_vector(31 downto 0);
    divisor:in std_logic_vector(7 downto 0);
    fractional:out std_logic_vector(7 downto 0);
    quotient:out std_logic_vector(31 downto 0);
    rfd:out std_logic
  );
end xldivider_generator_4c82698e6ec63d36ca8d57faf12d4ed2;


architecture behavior of xldivider_generator_4c82698e6ec63d36ca8d57faf12d4ed2  is
  component dv_gn_v3_0_56e83f20db65428d
    port(
      ce:in std_logic;
      clk:in std_logic;
      dividend:in std_logic_vector(31 downto 0);
      divisor:in std_logic_vector(7 downto 0);
      fractional:out std_logic_vector(7 downto 0);
      quotient:out std_logic_vector(31 downto 0);
      rfd:out std_logic
    );
end component;
begin
  dv_gn_v3_0_56e83f20db65428d_instance : dv_gn_v3_0_56e83f20db65428d
    port map(
      ce=>ce,
      clk=>clk,
      dividend=>dividend,
      divisor=>divisor,
      fractional=>fractional,
      quotient=>quotient,
      rfd=>rfd
    );
end  behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library thread_id_calc_lib;
use thread_id_calc_lib.conv_pkg.all;

entity xldivider_generator_2f6e135f81dffa050d9566043f612864 is 
  port(
    ce:in std_logic;
    clk:in std_logic;
    dividend:in std_logic_vector(5 downto 0);
    divisor:in std_logic_vector(7 downto 0);
    fractional:out std_logic_vector(7 downto 0);
    quotient:out std_logic_vector(5 downto 0);
    rfd:out std_logic
  );
end xldivider_generator_2f6e135f81dffa050d9566043f612864;


architecture behavior of xldivider_generator_2f6e135f81dffa050d9566043f612864  is
  component dv_gn_v3_0_26253f791d7c00ab
    port(
      ce:in std_logic;
      clk:in std_logic;
      dividend:in std_logic_vector(5 downto 0);
      divisor:in std_logic_vector(7 downto 0);
      fractional:out std_logic_vector(7 downto 0);
      quotient:out std_logic_vector(5 downto 0);
      rfd:out std_logic
    );
end component;
begin
  dv_gn_v3_0_26253f791d7c00ab_instance : dv_gn_v3_0_26253f791d7c00ab
    port map(
      ce=>ce,
      clk=>clk,
      dividend=>dividend,
      divisor=>divisor,
      fractional=>fractional,
      quotient=>quotient,
      rfd=>rfd
    );
end  behavior;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
library thread_id_calc_lib;
use thread_id_calc_lib.conv_pkg.all;

entity xldivider_generator_8dc90e2097a0b607ad0483b6293f4ad3 is 
  port(
    ce:in std_logic;
    clk:in std_logic;
    dividend:in std_logic_vector(31 downto 0);
    divisor:in std_logic_vector(5 downto 0);
    fractional:out std_logic_vector(5 downto 0);
    quotient:out std_logic_vector(31 downto 0);
    rfd:out std_logic
  );
end xldivider_generator_8dc90e2097a0b607ad0483b6293f4ad3;


architecture behavior of xldivider_generator_8dc90e2097a0b607ad0483b6293f4ad3  is
  component dv_gn_v3_0_90662698f61d80cb
    port(
      ce:in std_logic;
      clk:in std_logic;
      dividend:in std_logic_vector(31 downto 0);
      divisor:in std_logic_vector(5 downto 0);
      fractional:out std_logic_vector(5 downto 0);
      quotient:out std_logic_vector(31 downto 0);
      rfd:out std_logic
    );
end component;
begin
  dv_gn_v3_0_90662698f61d80cb_instance : dv_gn_v3_0_90662698f61d80cb
    port map(
      ce=>ce,
      clk=>clk,
      dividend=>dividend,
      divisor=>divisor,
      fractional=>fractional,
      quotient=>quotient,
      rfd=>rfd
    );
end  behavior;

library IEEE;
use IEEE.std_logic_1164.all;
library thread_id_calc_lib;
use thread_id_calc_lib.conv_pkg.all;

-- Generated from Simulink block "thread_id_calc"

entity thread_id_calc is
  port (
    block_indx_in: in std_logic_vector(15 downto 0); 
    block_x_in: in std_logic_vector(15 downto 0); 
    block_y_in: in std_logic_vector(15 downto 0); 
    block_z_in: in std_logic_vector(15 downto 0); 
    ce_1: in std_logic; 
    clk_1: in std_logic; 
    en: in std_logic; 
    num_cores_in: in std_logic_vector(7 downto 0); 
    warp_size_in: in std_logic_vector(5 downto 0); 
    warps_per_block_in: in std_logic_vector(5 downto 0); 
    x_indx_in: in std_logic_vector(15 downto 0); 
    y_indx_in: in std_logic_vector(15 downto 0); 
    z_indx_in: in std_logic_vector(15 downto 0); 
    data_valid: out std_logic; 
    thread_id_out: out std_logic_vector(31 downto 0); 
    thread_lane_id_out: out std_logic_vector(7 downto 0); 
    warp_id_out: out std_logic_vector(31 downto 0); 
    warp_lane_id_out: out std_logic_vector(5 downto 0)
  );
end thread_id_calc;

architecture structural of thread_id_calc is
  attribute core_generation_info: string;
  attribute core_generation_info of structural : architecture is "thread_id_calc,sysgen_core,{clock_period=10.00000000,clocking=Clock_Enables,compilation=NGC_Netlist,sample_periods=1.00000000000,testbench=1,total_blocks=66,xilinx_adder_subtracter_block=3,xilinx_arithmetic_relational_operator_block=1,xilinx_binary_shift_operator_block=2,xilinx_constant_block_block=1,xilinx_counter_block=1,xilinx_delay_block=1,xilinx_divider_generator_3_0_block=3,xilinx_gateway_in_block=11,xilinx_gateway_out_block=5,xilinx_logical_block_block=1,xilinx_multiplier_block=3,xilinx_register_block=15,xilinx_resource_estimator_block=1,xilinx_system_generator_block=1,xilinx_type_converter_block=1,}";

  signal addsub_s_net: std_logic_vector(31 downto 0);
  signal block_indx_in_net: std_logic_vector(15 downto 0);
  signal block_x_in_net: std_logic_vector(15 downto 0);
  signal block_y_in_net: std_logic_vector(15 downto 0);
  signal block_z_in_net: std_logic_vector(15 downto 0);
  signal ce_1_sg_x0: std_logic;
  signal clk_1_sg_x0: std_logic;
  signal constant_op_net: std_logic_vector(7 downto 0);
  signal convert_dout_net: std_logic;
  signal counter_op_net: std_logic_vector(7 downto 0);
  signal data_valid_net: std_logic;
  signal delay_q_net: std_logic_vector(21 downto 0);
  signal en_net: std_logic;
  signal lane_id_o1_quotient_net: std_logic_vector(5 downto 0);
  signal lane_id_o_fractional_net: std_logic_vector(7 downto 0);
  signal logical_y_net: std_logic_vector(31 downto 0);
  signal mult1_p_net: std_logic_vector(31 downto 0);
  signal mult2_p_net: std_logic_vector(21 downto 0);
  signal mult_p_net: std_logic_vector(31 downto 0);
  signal num_cores_in_net: std_logic_vector(7 downto 0);
  signal register10_q_net: std_logic_vector(7 downto 0);
  signal register1_q_net: std_logic_vector(15 downto 0);
  signal register2_q_net: std_logic_vector(15 downto 0);
  signal register3_q_net: std_logic_vector(15 downto 0);
  signal register4_q_net: std_logic_vector(15 downto 0);
  signal register5_q_net: std_logic_vector(15 downto 0);
  signal register7_q_net: std_logic_vector(5 downto 0);
  signal register8_q_net: std_logic_vector(5 downto 0);
  signal register9_q_net: std_logic;
  signal register_q_net: std_logic_vector(15 downto 0);
  signal shift1_op_net: std_logic_vector(31 downto 0);
  signal shift_op_net: std_logic_vector(31 downto 0);
  signal thread_id_o_s_net: std_logic_vector(31 downto 0);
  signal thread_id_out_net: std_logic_vector(31 downto 0);
  signal thread_lane_id_out_net: std_logic_vector(7 downto 0);
  signal warp_id_o1_fractional_net: std_logic_vector(5 downto 0);
  signal warp_id_o1_quotient_net: std_logic_vector(31 downto 0);
  signal warp_id_o_s_net: std_logic_vector(31 downto 0);
  signal warp_id_out_net: std_logic_vector(31 downto 0);
  signal warp_lane_id_out_net: std_logic_vector(5 downto 0);
  signal warp_size_in_net: std_logic_vector(5 downto 0);
  signal warps_per_block_in_net: std_logic_vector(5 downto 0);
  signal x_indx_in_net: std_logic_vector(15 downto 0);
  signal y_indx_in_net: std_logic_vector(15 downto 0);
  signal z_indx_in_net: std_logic_vector(15 downto 0);

begin
  block_indx_in_net <= block_indx_in;
  block_x_in_net <= block_x_in;
  block_y_in_net <= block_y_in;
  block_z_in_net <= block_z_in;
  ce_1_sg_x0 <= ce_1;
  clk_1_sg_x0 <= clk_1;
  en_net <= en;
  num_cores_in_net <= num_cores_in;
  warp_size_in_net <= warp_size_in;
  warps_per_block_in_net <= warps_per_block_in;
  x_indx_in_net <= x_indx_in;
  y_indx_in_net <= y_indx_in;
  z_indx_in_net <= z_indx_in;
  data_valid <= data_valid_net;
  thread_id_out <= thread_id_out_net;
  thread_lane_id_out <= thread_lane_id_out_net;
  warp_id_out <= warp_id_out_net;
  warp_lane_id_out <= warp_lane_id_out_net;

  addsub: entity thread_id_calc_lib.xladdsub
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 16,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 32,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 33,
      core_name0 => "addsb_11_0_f45daeb7eb283db0",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 33,
      latency => 0,
      overflow => 2,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 32
    )
    port map (
      a => register1_q_net,
      b => mult_p_net,
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      en => "1",
      s => addsub_s_net
    );

  constant_x0: entity thread_id_calc_lib.constant_7db069ad14
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      op => constant_op_net
    );

  convert: entity thread_id_calc_lib.xlconvert
    generic map (
      bool_conversion => 1,
      din_arith => 1,
      din_bin_pt => 0,
      din_width => 1,
      dout_arith => 1,
      dout_bin_pt => 0,
      dout_width => 1,
      latency => 0,
      overflow => xlWrap,
      quantization => xlTruncate
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      din(0) => en_net,
      en => "1",
      dout(0) => convert_dout_net
    );

  counter: entity thread_id_calc_lib.xlcounter_free
    generic map (
      core_name0 => "cntr_11_0_e7514e290b172ea1",
      op_arith => xlUnsigned,
      op_width => 8
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      en(0) => register9_q_net,
      rst(0) => data_valid_net,
      op => counter_op_net
    );

  delay: entity thread_id_calc_lib.xldelay
    generic map (
      latency => 3,
      reg_retiming => 0,
      width => 22
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d => mult2_p_net,
      en => '1',
      q => delay_q_net
    );

  lane_id_o: entity thread_id_calc_lib.xldivider_generator_4c82698e6ec63d36ca8d57faf12d4ed2
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      dividend => thread_id_o_s_net,
      divisor => register10_q_net,
      fractional => lane_id_o_fractional_net
    );

  lane_id_o1: entity thread_id_calc_lib.xldivider_generator_2f6e135f81dffa050d9566043f612864
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      dividend => warp_id_o1_fractional_net,
      divisor => register10_q_net,
      quotient => lane_id_o1_quotient_net
    );

  logical: entity thread_id_calc_lib.logical_0d8e48dd8a
    port map (
      ce => '0',
      clk => '0',
      clr => '0',
      d0 => register_q_net,
      d1 => shift1_op_net,
      d2 => shift_op_net,
      y => logical_y_net
    );

  mult: entity thread_id_calc_lib.xlmult
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 16,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 16,
      c_a_type => 1,
      c_a_width => 16,
      c_b_type => 1,
      c_b_width => 16,
      c_baat => 16,
      c_output_width => 32,
      c_type => 1,
      core_name0 => "mult_11_2_7165ba8b8713bab6",
      extra_registers => 0,
      multsign => 1,
      overflow => 2,
      p_arith => xlUnsigned,
      p_bin_pt => 0,
      p_width => 32,
      quantization => 1
    )
    port map (
      a => register2_q_net,
      b => register5_q_net,
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      core_ce => ce_1_sg_x0,
      core_clk => clk_1_sg_x0,
      core_clr => '1',
      en => "1",
      rst => "0",
      p => mult_p_net
    );

  mult1: entity thread_id_calc_lib.xlmult
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 32,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 16,
      c_a_type => 1,
      c_a_width => 32,
      c_b_type => 1,
      c_b_width => 16,
      c_baat => 32,
      c_output_width => 48,
      c_type => 1,
      core_name0 => "mult_11_2_3f458b247f28c718",
      extra_registers => 1,
      multsign => 1,
      overflow => 2,
      p_arith => xlUnsigned,
      p_bin_pt => 0,
      p_width => 32,
      quantization => 1
    )
    port map (
      a => addsub_s_net,
      b => register4_q_net,
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      core_ce => ce_1_sg_x0,
      core_clk => clk_1_sg_x0,
      core_clr => '1',
      en => "1",
      rst => "0",
      p => mult1_p_net
    );

  mult2: entity thread_id_calc_lib.xlmult
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 16,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 6,
      c_a_type => 1,
      c_a_width => 16,
      c_b_type => 1,
      c_b_width => 6,
      c_baat => 16,
      c_output_width => 22,
      c_type => 1,
      core_name0 => "mult_11_2_234eb26fa92ee3d2",
      extra_registers => 0,
      multsign => 1,
      overflow => 1,
      p_arith => xlUnsigned,
      p_bin_pt => 0,
      p_width => 22,
      quantization => 1
    )
    port map (
      a => register3_q_net,
      b => register8_q_net,
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      core_ce => ce_1_sg_x0,
      core_clk => clk_1_sg_x0,
      core_clr => '1',
      en => "1",
      rst => "0",
      p => mult2_p_net
    );

  register1: entity thread_id_calc_lib.xlregister
    generic map (
      d_width => 16,
      init_value => b"0000000000000000"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d => y_indx_in_net,
      en(0) => convert_dout_net,
      rst => "0",
      q => register1_q_net
    );

  register10: entity thread_id_calc_lib.xlregister
    generic map (
      d_width => 8,
      init_value => b"00000000"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d => num_cores_in_net,
      en(0) => convert_dout_net,
      rst => "0",
      q => register10_q_net
    );

  register11: entity thread_id_calc_lib.xlregister
    generic map (
      d_width => 32,
      init_value => b"00000000000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d => logical_y_net,
      en(0) => data_valid_net,
      rst => "0",
      q => thread_id_out_net
    );

  register12: entity thread_id_calc_lib.xlregister
    generic map (
      d_width => 32,
      init_value => b"00000000000000000000000000000000"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d => warp_id_o_s_net,
      en(0) => data_valid_net,
      rst => "0",
      q => warp_id_out_net
    );

  register13: entity thread_id_calc_lib.xlregister
    generic map (
      d_width => 6,
      init_value => b"000000"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d => lane_id_o1_quotient_net,
      en(0) => data_valid_net,
      rst => "0",
      q => warp_lane_id_out_net
    );

  register14: entity thread_id_calc_lib.xlregister
    generic map (
      d_width => 8,
      init_value => b"00000000"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d => lane_id_o_fractional_net,
      en(0) => data_valid_net,
      rst => "0",
      q => thread_lane_id_out_net
    );

  register2: entity thread_id_calc_lib.xlregister
    generic map (
      d_width => 16,
      init_value => b"0000000000000000"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d => z_indx_in_net,
      en(0) => convert_dout_net,
      rst => "0",
      q => register2_q_net
    );

  register3: entity thread_id_calc_lib.xlregister
    generic map (
      d_width => 16,
      init_value => b"0000000000000000"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d => block_indx_in_net,
      en(0) => convert_dout_net,
      rst => "0",
      q => register3_q_net
    );

  register4: entity thread_id_calc_lib.xlregister
    generic map (
      d_width => 16,
      init_value => b"0000000000000000"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d => block_x_in_net,
      en(0) => convert_dout_net,
      rst => "0",
      q => register4_q_net
    );

  register5: entity thread_id_calc_lib.xlregister
    generic map (
      d_width => 16,
      init_value => b"0000000000000000"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d => block_y_in_net,
      en(0) => convert_dout_net,
      rst => "0",
      q => register5_q_net
    );

  register7: entity thread_id_calc_lib.xlregister
    generic map (
      d_width => 6,
      init_value => b"000000"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d => warp_size_in_net,
      en(0) => convert_dout_net,
      rst => "0",
      q => register7_q_net
    );

  register8: entity thread_id_calc_lib.xlregister
    generic map (
      d_width => 6,
      init_value => b"000000"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d => warps_per_block_in_net,
      en(0) => convert_dout_net,
      rst => "0",
      q => register8_q_net
    );

  register9: entity thread_id_calc_lib.xlregister
    generic map (
      d_width => 1,
      init_value => b"0"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d(0) => convert_dout_net,
      en(0) => convert_dout_net,
      rst(0) => data_valid_net,
      q(0) => register9_q_net
    );

  register_x0: entity thread_id_calc_lib.xlregister
    generic map (
      d_width => 16,
      init_value => b"0000000000000000"
    )
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      d => x_indx_in_net,
      en(0) => convert_dout_net,
      rst => "0",
      q => register_q_net
    );

  relational: entity thread_id_calc_lib.relational_54048c8b02
    port map (
      a => counter_op_net,
      b => constant_op_net,
      ce => '0',
      clk => '0',
      clr => '0',
      op(0) => data_valid_net
    );

  shift: entity thread_id_calc_lib.shift_63b52ec892
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      ip => register2_q_net,
      op => shift_op_net
    );

  shift1: entity thread_id_calc_lib.shift_cdf6c3fa1e
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      ip => register1_q_net,
      op => shift1_op_net
    );

  thread_id_o: entity thread_id_calc_lib.xladdsub
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 16,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 32,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 33,
      core_name0 => "addsb_11_0_f45daeb7eb283db0",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 33,
      latency => 0,
      overflow => 2,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 32
    )
    port map (
      a => register_q_net,
      b => mult1_p_net,
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      en => "1",
      s => thread_id_o_s_net
    );

  warp_id_o: entity thread_id_calc_lib.xladdsub
    generic map (
      a_arith => xlUnsigned,
      a_bin_pt => 0,
      a_width => 32,
      b_arith => xlUnsigned,
      b_bin_pt => 0,
      b_width => 22,
      c_has_c_out => 0,
      c_latency => 0,
      c_output_width => 33,
      core_name0 => "addsb_11_0_f45daeb7eb283db0",
      extra_registers => 0,
      full_s_arith => 1,
      full_s_width => 33,
      latency => 0,
      overflow => 2,
      quantization => 1,
      s_arith => xlUnsigned,
      s_bin_pt => 0,
      s_width => 32
    )
    port map (
      a => warp_id_o1_quotient_net,
      b => delay_q_net,
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      clr => '0',
      en => "1",
      s => warp_id_o_s_net
    );

  warp_id_o1: entity thread_id_calc_lib.xldivider_generator_8dc90e2097a0b607ad0483b6293f4ad3
    port map (
      ce => ce_1_sg_x0,
      clk => clk_1_sg_x0,
      dividend => thread_id_o_s_net,
      divisor => register7_q_net,
      fractional => warp_id_o1_fractional_net,
      quotient => warp_id_o1_quotient_net
    );

end structural;
